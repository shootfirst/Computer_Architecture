module IF(
  input         clock,
  input         reset,
  output [31:0] io_mmu_addr,
  output [3:0]  io_mmu_mode,
  input  [31:0] io_mmu_rdata,
  input         io_mmu_ok,
  input         io_mmu_pageFault,
  output [31:0] io_id_inst,
  output        io_id_excep_valid,
  output [31:0] io_id_excep_code,
  output [31:0] io_id_excep_value,
  output [31:0] io_id_excep_pc,
  output        io_id_excep_valid_inst,
  input         io_id_branch_valid,
  input  [31:0] io_id_branch_bits,
  input         io_id_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[IF.scala 13:27]
  reg  log_branch_valid; // @[IF.scala 14:27]
  reg [31:0] log_branch_bits; // @[IF.scala 14:27]
  reg  log_inst_valid; // @[IF.scala 15:27]
  reg [31:0] log_inst_bits; // @[IF.scala 15:27]
  wire  branch_valid = io_id_branch_valid ? io_id_branch_valid : log_branch_valid; // @[IF.scala 21:19]
  wire  inst_valid = log_inst_valid ? log_inst_valid : io_mmu_ok; // @[IF.scala 22:19]
  wire [31:0] inst_bits = log_inst_valid ? log_inst_bits : io_mmu_rdata; // @[IF.scala 22:19]
  wire  _T_2 = ~log_inst_valid; // @[IF.scala 28:8]
  wire  _T_3 = _T_2 & io_mmu_ok; // @[IF.scala 28:24]
  wire  _GEN_2 = _T_3 | log_inst_valid; // @[IF.scala 28:38]
  wire  _T_4 = ~inst_valid; // @[IF.scala 33:15]
  wire  _T_5 = ~io_id_ready; // @[IF.scala 33:30]
  wire  stall = _T_4 | _T_5; // @[IF.scala 33:27]
  wire  _T_6 = ~stall; // @[IF.scala 36:8]
  wire [31:0] _T_8 = pc + 32'h4; // @[IF.scala 39:25]
  wire  _T_12 = log_inst_valid ? 1'h0 : 1'h1; // @[IF.scala 46:22]
  wire  _T_14 = stall | branch_valid; // @[IF.scala 55:16]
  wire  _T_15 = ~_T_14; // @[IF.scala 55:8]
  wire  _T_17 = |pc[1:0]; // @[IF.scala 59:18]
  wire [31:0] _GEN_10 = _T_17 ? pc : 32'h0; // @[IF.scala 59:23]
  wire  _GEN_12 = io_mmu_pageFault | _T_17; // @[IF.scala 64:28]
  wire [31:0] _GEN_13 = io_mmu_pageFault ? pc : _GEN_10; // @[IF.scala 64:28]
  wire [31:0] _GEN_14 = io_mmu_pageFault ? 32'hc : 32'h0; // @[IF.scala 64:28]
  assign io_mmu_addr = pc; // @[IF.scala 45:16]
  assign io_mmu_mode = {{3'd0}, _T_12}; // @[IF.scala 46:16]
  assign io_id_inst = _T_15 ? inst_bits : 32'h13; // @[IF.scala 52:15 IF.scala 56:16]
  assign io_id_excep_valid = _T_15 & _GEN_12; // @[IF.scala 53:15 IF.scala 60:25 IF.scala 65:25]
  assign io_id_excep_code = _T_15 ? _GEN_14 : 32'h0; // @[IF.scala 53:15 IF.scala 62:24 IF.scala 67:24]
  assign io_id_excep_value = _T_15 ? _GEN_13 : 32'h0; // @[IF.scala 53:15 IF.scala 61:25 IF.scala 66:25]
  assign io_id_excep_pc = _T_15 ? pc : 32'h0; // @[IF.scala 53:15 IF.scala 57:20]
  assign io_id_excep_valid_inst = ~_T_14; // @[IF.scala 53:15 IF.scala 58:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  log_branch_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  log_branch_bits = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  log_inst_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  log_inst_bits = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h80000000;
    end else if (_T_6) begin
      if (branch_valid) begin
        if (io_id_branch_valid) begin
          pc <= io_id_branch_bits;
        end else begin
          pc <= log_branch_bits;
        end
      end else begin
        pc <= _T_8;
      end
    end
    if (reset) begin
      log_branch_valid <= 1'h0;
    end else if (_T_6) begin
      log_branch_valid <= 1'h0;
    end else if (io_id_branch_valid) begin
      log_branch_valid <= io_id_branch_valid;
    end
    if (reset) begin
      log_branch_bits <= 32'h0;
    end else if (_T_6) begin
      log_branch_bits <= 32'h0;
    end else if (io_id_branch_valid) begin
      log_branch_bits <= io_id_branch_bits;
    end
    if (reset) begin
      log_inst_valid <= 1'h0;
    end else if (_T_6) begin
      log_inst_valid <= 1'h0;
    end else begin
      log_inst_valid <= _GEN_2;
    end
    if (reset) begin
      log_inst_bits <= 32'h0;
    end else if (_T_6) begin
      log_inst_bits <= 32'h0;
    end else if (_T_3) begin
      log_inst_bits <= io_mmu_rdata;
    end
  end
endmodule
module ID(
  input         clock,
  input         reset,
  input  [31:0] io_iff_inst,
  input         io_iff_excep_valid,
  input  [31:0] io_iff_excep_code,
  input  [31:0] io_iff_excep_value,
  input  [31:0] io_iff_excep_pc,
  input         io_iff_excep_valid_inst,
  output        io_iff_branch_valid,
  output [31:0] io_iff_branch_bits,
  output        io_iff_ready,
  output [4:0]  io_reg_read1_addr,
  input  [31:0] io_reg_read1_data,
  output [4:0]  io_reg_read2_addr,
  input  [31:0] io_reg_read2_data,
  output [31:0] io_ex_aluOp_rd1,
  output [31:0] io_ex_aluOp_rd2,
  output [4:0]  io_ex_aluOp_opt,
  output [4:0]  io_ex_wrRegOp_addr,
  output        io_ex_wrCSROp_valid,
  output [11:0] io_ex_wrCSROp_addr,
  output [31:0] io_ex_wrCSROp_data,
  output [31:0] io_ex_store_data,
  output        io_ex_excep_valid,
  output [31:0] io_ex_excep_code,
  output [31:0] io_ex_excep_value,
  output [31:0] io_ex_excep_pc,
  output        io_ex_excep_valid_inst,
  input         io_ex_ready,
  output [11:0] io_csr_addr,
  input  [31:0] io_csr_rdata,
  input  [1:0]  io_csr_prv,
  input         io_flush,
  input  [4:0]  io_exWrRegOp_addr,
  input  [31:0] io_exWrRegOp_data,
  input         io_exWrRegOp_rdy,
  input  [4:0]  io_memWrRegOp_addr,
  input  [31:0] io_memWrRegOp_data,
  input         io_exWrCSROp_valid,
  input  [11:0] io_exWrCSROp_addr,
  input  [31:0] io_exWrCSROp_data,
  input         io_memWrCSROp_valid,
  input  [11:0] io_memWrCSROp_addr,
  input  [31:0] io_memWrCSROp_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] inst; // @[ID.scala 37:22]
  reg  excep_valid; // @[ID.scala 38:22]
  reg [31:0] excep_code; // @[ID.scala 38:22]
  reg [31:0] excep_value; // @[ID.scala 38:22]
  reg [31:0] excep_pc; // @[ID.scala 38:22]
  reg  excep_valid_inst; // @[ID.scala 38:22]
  reg [1:0] fenceICnt; // @[ID.scala 40:26]
  wire  _T_223 = ~io_exWrRegOp_rdy; // @[ID.scala 122:13]
  wire  _T_224 = |io_exWrRegOp_addr; // @[ID.scala 122:54]
  wire  _T_225 = _T_223 & _T_224; // @[ID.scala 122:32]
  wire [4:0] rs1Addr = inst[19:15]; // @[ID.scala 65:22]
  wire  _T_209 = rs1Addr == io_exWrRegOp_addr; // @[ID.scala 118:28]
  wire [31:0] _T_2 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 32'h13 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 32'h2013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_7 = 32'h3013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_9 = 32'h4013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_11 = 32'h6013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 32'h7013 == _T_2; // @[Lookup.scala 31:38]
  wire [31:0] _T_14 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_15 = 32'h1013 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_17 = 32'h5013 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_19 = 32'h40005013 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_21 = 32'h33 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_23 = 32'h40000033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_25 = 32'h1033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_27 = 32'h2033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_29 = 32'h3033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_31 = 32'h4033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_33 = 32'h5033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h40005033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h6033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h7033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h3 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h1003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h2003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h4003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h5003 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h23 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h1023 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h2023 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h63 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h1063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h4063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h5063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h6063 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h7063 == _T_2; // @[Lookup.scala 31:38]
  wire [31:0] _T_68 = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h37 == _T_68; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h17 == _T_68; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h6f == _T_68; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'h67 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h73 == _T_68; // @[Lookup.scala 31:38]
  wire [31:0] _T_78 = inst & 32'hf00fffff; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'hf == _T_78; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h100f == inst; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'h2000033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'h2001033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h2002033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h2004033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h2005033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h2006033 == _T_14; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'h2007033 == _T_14; // @[Lookup.scala 31:38]
  wire [3:0] _T_96 = _T_95 ? 4'h1 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_97 = _T_93 ? 4'h1 : _T_96; // @[Lookup.scala 33:37]
  wire [3:0] _T_98 = _T_91 ? 4'h1 : _T_97; // @[Lookup.scala 33:37]
  wire [3:0] _T_99 = _T_89 ? 4'h1 : _T_98; // @[Lookup.scala 33:37]
  wire [3:0] _T_100 = _T_87 ? 4'h1 : _T_99; // @[Lookup.scala 33:37]
  wire [3:0] _T_101 = _T_85 ? 4'h1 : _T_100; // @[Lookup.scala 33:37]
  wire [3:0] _T_102 = _T_83 ? 4'h1 : _T_101; // @[Lookup.scala 33:37]
  wire [3:0] _T_103 = _T_81 ? 4'h8 : _T_102; // @[Lookup.scala 33:37]
  wire [3:0] _T_104 = _T_79 ? 4'h8 : _T_103; // @[Lookup.scala 33:37]
  wire [3:0] _T_105 = _T_77 ? 4'h7 : _T_104; // @[Lookup.scala 33:37]
  wire [3:0] _T_106 = _T_75 ? 4'h2 : _T_105; // @[Lookup.scala 33:37]
  wire [3:0] _T_107 = _T_73 ? 4'h6 : _T_106; // @[Lookup.scala 33:37]
  wire [3:0] _T_108 = _T_71 ? 4'h5 : _T_107; // @[Lookup.scala 33:37]
  wire [3:0] _T_109 = _T_69 ? 4'h5 : _T_108; // @[Lookup.scala 33:37]
  wire [3:0] _T_110 = _T_67 ? 4'h4 : _T_109; // @[Lookup.scala 33:37]
  wire [3:0] _T_111 = _T_65 ? 4'h4 : _T_110; // @[Lookup.scala 33:37]
  wire [3:0] _T_112 = _T_63 ? 4'h4 : _T_111; // @[Lookup.scala 33:37]
  wire [3:0] _T_113 = _T_61 ? 4'h4 : _T_112; // @[Lookup.scala 33:37]
  wire [3:0] _T_114 = _T_59 ? 4'h4 : _T_113; // @[Lookup.scala 33:37]
  wire [3:0] _T_115 = _T_57 ? 4'h4 : _T_114; // @[Lookup.scala 33:37]
  wire [3:0] _T_116 = _T_55 ? 4'h3 : _T_115; // @[Lookup.scala 33:37]
  wire [3:0] _T_117 = _T_53 ? 4'h3 : _T_116; // @[Lookup.scala 33:37]
  wire [3:0] _T_118 = _T_51 ? 4'h3 : _T_117; // @[Lookup.scala 33:37]
  wire [3:0] _T_119 = _T_49 ? 4'h2 : _T_118; // @[Lookup.scala 33:37]
  wire [3:0] _T_120 = _T_47 ? 4'h2 : _T_119; // @[Lookup.scala 33:37]
  wire [3:0] _T_121 = _T_45 ? 4'h2 : _T_120; // @[Lookup.scala 33:37]
  wire [3:0] _T_122 = _T_43 ? 4'h2 : _T_121; // @[Lookup.scala 33:37]
  wire [3:0] _T_123 = _T_41 ? 4'h2 : _T_122; // @[Lookup.scala 33:37]
  wire [3:0] _T_124 = _T_39 ? 4'h1 : _T_123; // @[Lookup.scala 33:37]
  wire [3:0] _T_125 = _T_37 ? 4'h1 : _T_124; // @[Lookup.scala 33:37]
  wire [3:0] _T_126 = _T_35 ? 4'h1 : _T_125; // @[Lookup.scala 33:37]
  wire [3:0] _T_127 = _T_33 ? 4'h1 : _T_126; // @[Lookup.scala 33:37]
  wire [3:0] _T_128 = _T_31 ? 4'h1 : _T_127; // @[Lookup.scala 33:37]
  wire [3:0] _T_129 = _T_29 ? 4'h1 : _T_128; // @[Lookup.scala 33:37]
  wire [3:0] _T_130 = _T_27 ? 4'h1 : _T_129; // @[Lookup.scala 33:37]
  wire [3:0] _T_131 = _T_25 ? 4'h1 : _T_130; // @[Lookup.scala 33:37]
  wire [3:0] _T_132 = _T_23 ? 4'h1 : _T_131; // @[Lookup.scala 33:37]
  wire [3:0] _T_133 = _T_21 ? 4'h1 : _T_132; // @[Lookup.scala 33:37]
  wire [3:0] _T_134 = _T_19 ? 4'h2 : _T_133; // @[Lookup.scala 33:37]
  wire [3:0] _T_135 = _T_17 ? 4'h2 : _T_134; // @[Lookup.scala 33:37]
  wire [3:0] _T_136 = _T_15 ? 4'h2 : _T_135; // @[Lookup.scala 33:37]
  wire [3:0] _T_137 = _T_13 ? 4'h2 : _T_136; // @[Lookup.scala 33:37]
  wire [3:0] _T_138 = _T_11 ? 4'h2 : _T_137; // @[Lookup.scala 33:37]
  wire [3:0] _T_139 = _T_9 ? 4'h2 : _T_138; // @[Lookup.scala 33:37]
  wire [3:0] _T_140 = _T_7 ? 4'h2 : _T_139; // @[Lookup.scala 33:37]
  wire [3:0] _T_141 = _T_5 ? 4'h2 : _T_140; // @[Lookup.scala 33:37]
  wire [3:0] decRes_0 = _T_3 ? 4'h2 : _T_141; // @[Lookup.scala 33:37]
  wire  _T_210 = 4'h1 == decRes_0; // @[ID.scala 119:34]
  wire  _T_211 = 4'h2 == decRes_0; // @[ID.scala 119:34]
  wire  _T_214 = _T_210 | _T_211; // @[ID.scala 119:57]
  wire  _T_212 = 4'h3 == decRes_0; // @[ID.scala 119:34]
  wire  _T_215 = _T_214 | _T_212; // @[ID.scala 119:57]
  wire  _T_213 = 4'h4 == decRes_0; // @[ID.scala 119:34]
  wire  _T_216 = _T_215 | _T_213; // @[ID.scala 119:57]
  wire  rs1Hazard = _T_209 & _T_216; // @[ID.scala 118:51]
  wire [4:0] rs2Addr = inst[24:20]; // @[ID.scala 66:22]
  wire  _T_217 = rs2Addr == io_exWrRegOp_addr; // @[ID.scala 120:28]
  wire  _T_221 = _T_210 | _T_212; // @[ID.scala 121:57]
  wire  _T_222 = _T_221 | _T_213; // @[ID.scala 121:57]
  wire  rs2Hazard = _T_217 & _T_222; // @[ID.scala 120:51]
  wire  _T_226 = rs1Hazard | rs2Hazard; // @[ID.scala 122:73]
  wire  _T_227 = _T_225 & _T_226; // @[ID.scala 122:59]
  wire  _T_228 = ~io_ex_ready; // @[ID.scala 122:90]
  wire  stall = _T_227 | _T_228; // @[ID.scala 122:87]
  wire [4:0] _T_142 = _T_95 ? 5'h12 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_143 = _T_93 ? 5'h11 : _T_142; // @[Lookup.scala 33:37]
  wire [4:0] _T_144 = _T_91 ? 5'h10 : _T_143; // @[Lookup.scala 33:37]
  wire [4:0] _T_145 = _T_89 ? 5'hf : _T_144; // @[Lookup.scala 33:37]
  wire [4:0] _T_146 = _T_87 ? 5'hd : _T_145; // @[Lookup.scala 33:37]
  wire [4:0] _T_147 = _T_85 ? 5'hc : _T_146; // @[Lookup.scala 33:37]
  wire [4:0] _T_148 = _T_83 ? 5'hb : _T_147; // @[Lookup.scala 33:37]
  wire [4:0] _T_149 = _T_81 ? 5'h0 : _T_148; // @[Lookup.scala 33:37]
  wire [4:0] _T_150 = _T_79 ? 5'h0 : _T_149; // @[Lookup.scala 33:37]
  wire [4:0] _T_151 = _T_77 ? 5'h0 : _T_150; // @[Lookup.scala 33:37]
  wire [4:0] _T_152 = _T_75 ? 5'ha : _T_151; // @[Lookup.scala 33:37]
  wire [4:0] _T_153 = _T_73 ? 5'h0 : _T_152; // @[Lookup.scala 33:37]
  wire [4:0] _T_154 = _T_71 ? 5'h1 : _T_153; // @[Lookup.scala 33:37]
  wire [4:0] _T_155 = _T_69 ? 5'h0 : _T_154; // @[Lookup.scala 33:37]
  wire [4:0] _T_156 = _T_67 ? 5'h7 : _T_155; // @[Lookup.scala 33:37]
  wire [4:0] _T_157 = _T_65 ? 5'h9 : _T_156; // @[Lookup.scala 33:37]
  wire [4:0] _T_158 = _T_63 ? 5'h6 : _T_157; // @[Lookup.scala 33:37]
  wire [4:0] _T_159 = _T_61 ? 5'h8 : _T_158; // @[Lookup.scala 33:37]
  wire [4:0] _T_160 = _T_59 ? 5'ha : _T_159; // @[Lookup.scala 33:37]
  wire [4:0] _T_161 = _T_57 ? 5'h4 : _T_160; // @[Lookup.scala 33:37]
  wire [4:0] _T_162 = _T_55 ? 5'h14 : _T_161; // @[Lookup.scala 33:37]
  wire [4:0] _T_163 = _T_53 ? 5'h15 : _T_162; // @[Lookup.scala 33:37]
  wire [4:0] _T_164 = _T_51 ? 5'h16 : _T_163; // @[Lookup.scala 33:37]
  wire [4:0] _T_165 = _T_49 ? 5'h1b : _T_164; // @[Lookup.scala 33:37]
  wire [4:0] _T_166 = _T_47 ? 5'h1d : _T_165; // @[Lookup.scala 33:37]
  wire [4:0] _T_167 = _T_45 ? 5'h18 : _T_166; // @[Lookup.scala 33:37]
  wire [4:0] _T_168 = _T_43 ? 5'h1a : _T_167; // @[Lookup.scala 33:37]
  wire [4:0] _T_169 = _T_41 ? 5'h1c : _T_168; // @[Lookup.scala 33:37]
  wire [4:0] _T_170 = _T_39 ? 5'h6 : _T_169; // @[Lookup.scala 33:37]
  wire [4:0] _T_171 = _T_37 ? 5'h5 : _T_170; // @[Lookup.scala 33:37]
  wire [4:0] _T_172 = _T_35 ? 5'h9 : _T_171; // @[Lookup.scala 33:37]
  wire [4:0] _T_173 = _T_33 ? 5'h8 : _T_172; // @[Lookup.scala 33:37]
  wire [4:0] _T_174 = _T_31 ? 5'h4 : _T_173; // @[Lookup.scala 33:37]
  wire [4:0] _T_175 = _T_29 ? 5'h3 : _T_174; // @[Lookup.scala 33:37]
  wire [4:0] _T_176 = _T_27 ? 5'h2 : _T_175; // @[Lookup.scala 33:37]
  wire [4:0] _T_177 = _T_25 ? 5'h7 : _T_176; // @[Lookup.scala 33:37]
  wire [4:0] _T_178 = _T_23 ? 5'h1 : _T_177; // @[Lookup.scala 33:37]
  wire [4:0] _T_179 = _T_21 ? 5'h0 : _T_178; // @[Lookup.scala 33:37]
  wire [4:0] _T_180 = _T_19 ? 5'h9 : _T_179; // @[Lookup.scala 33:37]
  wire [4:0] _T_181 = _T_17 ? 5'h8 : _T_180; // @[Lookup.scala 33:37]
  wire [4:0] _T_182 = _T_15 ? 5'h7 : _T_181; // @[Lookup.scala 33:37]
  wire [4:0] _T_183 = _T_13 ? 5'h6 : _T_182; // @[Lookup.scala 33:37]
  wire [4:0] _T_184 = _T_11 ? 5'h5 : _T_183; // @[Lookup.scala 33:37]
  wire [4:0] _T_185 = _T_9 ? 5'h4 : _T_184; // @[Lookup.scala 33:37]
  wire [4:0] _T_186 = _T_7 ? 5'h3 : _T_185; // @[Lookup.scala 33:37]
  wire [4:0] _T_187 = _T_5 ? 5'h2 : _T_186; // @[Lookup.scala 33:37]
  wire [4:0] decRes_1 = _T_3 ? 5'h0 : _T_187; // @[Lookup.scala 33:37]
  wire [4:0] rdAddr = inst[11:7]; // @[ID.scala 67:22]
  wire [11:0] csrAddr = inst[31:20]; // @[ID.scala 68:22]
  wire  _T_188 = rs1Addr == 5'h0; // @[ID.scala 78:14]
  wire  _T_190 = rs1Addr == io_memWrRegOp_addr; // @[ID.scala 80:14]
  wire [31:0] _T_191 = _T_190 ? io_memWrRegOp_data : io_reg_read1_data; // @[Mux.scala 47:69]
  wire [31:0] _T_192 = _T_209 ? io_exWrRegOp_data : _T_191; // @[Mux.scala 47:69]
  wire [31:0] rs1Val = _T_188 ? 32'h0 : _T_192; // @[Mux.scala 47:69]
  wire  _T_193 = rs2Addr == 5'h0; // @[ID.scala 83:14]
  wire  _T_195 = rs2Addr == io_memWrRegOp_addr; // @[ID.scala 85:14]
  wire [31:0] _T_196 = _T_195 ? io_memWrRegOp_data : io_reg_read2_data; // @[Mux.scala 47:69]
  wire [31:0] _T_197 = _T_217 ? io_exWrRegOp_data : _T_196; // @[Mux.scala 47:69]
  wire [31:0] rs2Val = _T_193 ? 32'h0 : _T_197; // @[Mux.scala 47:69]
  wire  _T_198 = csrAddr == io_exWrCSROp_addr; // @[ID.scala 88:14]
  wire  _T_199 = _T_198 & io_exWrCSROp_valid; // @[ID.scala 88:36]
  wire  _T_200 = csrAddr == io_memWrCSROp_addr; // @[ID.scala 89:14]
  wire  _T_201 = _T_200 & io_memWrCSROp_valid; // @[ID.scala 89:37]
  wire [31:0] _T_202 = _T_201 ? io_memWrCSROp_data : io_csr_rdata; // @[Mux.scala 47:69]
  wire [31:0] csrVal = _T_199 ? io_exWrCSROp_data : _T_202; // @[Mux.scala 47:69]
  wire  _T_207 = ~stall; // @[ID.scala 108:49]
  wire [11:0] _T_233 = inst[31:20]; // @[ID.scala 155:28]
  wire [11:0] _T_248 = {inst[31:25],rdAddr}; // @[ID.scala 168:45]
  wire [12:0] _T_280 = {inst[31],inst[7],inst[30:25],inst[11:8],1'h0}; // @[ID.scala 180:75]
  wire  _T_287 = 4'h5 == decRes_0; // @[Conditional.scala 37:30]
  wire [31:0] _T_289 = inst & 32'hfffff000; // @[ID.scala 189:40]
  wire  _T_293 = 4'h6 == decRes_0; // @[Conditional.scala 37:30]
  wire [20:0] _T_302 = {inst[31],inst[19:12],inst[20],inst[30:21],1'h0}; // @[ID.scala 197:76]
  wire [20:0] _GEN_100 = _T_293 ? $signed(_T_302) : $signed(21'sh0); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_114 = _T_287 ? $signed(_T_289) : $signed({{11{_GEN_100[20]}},_GEN_100}); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_128 = _T_213 ? $signed({{19{_T_280[12]}},_T_280}) : $signed(_GEN_114); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_144 = _T_212 ? $signed({{20{_T_248[11]}},_T_248}) : $signed(_GEN_128); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_161 = _T_211 ? $signed({{20{_T_233[11]}},_T_233}) : $signed(_GEN_144); // @[Conditional.scala 39:67]
  wire [31:0] _GEN_181 = _T_210 ? $signed(32'sh0) : $signed(_GEN_161); // @[Conditional.scala 40:58]
  wire [31:0] _T_234 = stall ? $signed(32'sh0) : $signed(_GEN_181); // @[ID.scala 157:32]
  wire  _T_235 = decRes_1 == 5'ha; // @[ID.scala 160:35]
  wire [31:0] _T_238 = _T_234 + rs1Val; // @[ID.scala 161:36]
  wire [31:0] _T_240 = _T_238 & 32'hfffffffe; // @[ID.scala 161:46]
  wire  _T_242 = |_T_240[1:0]; // @[ID.scala 127:22]
  wire  _T_243 = ~excep_valid; // @[ID.scala 128:12]
  wire  _GEN_12 = _T_243 | excep_valid; // @[ID.scala 128:26]
  wire [31:0] _GEN_13 = _T_243 ? _T_240 : excep_value; // @[ID.scala 128:26]
  wire [31:0] _GEN_14 = _T_243 ? 32'h0 : excep_code; // @[ID.scala 128:26]
  wire  _GEN_15 = _T_242 ? _GEN_12 : excep_valid; // @[ID.scala 127:27]
  wire [31:0] _GEN_16 = _T_242 ? _GEN_13 : excep_value; // @[ID.scala 127:27]
  wire [31:0] _GEN_17 = _T_242 ? _GEN_14 : excep_code; // @[ID.scala 127:27]
  wire [31:0] _GEN_18 = _T_242 ? 32'h0 : _T_240; // @[ID.scala 127:27]
  wire  _GEN_19 = _T_242 ? 1'h0 : 1'h1; // @[ID.scala 127:27]
  wire  _GEN_20 = _T_235 ? _GEN_15 : excep_valid; // @[ID.scala 160:53]
  wire [31:0] _GEN_21 = _T_235 ? _GEN_16 : excep_value; // @[ID.scala 160:53]
  wire [31:0] _GEN_22 = _T_235 ? _GEN_17 : excep_code; // @[ID.scala 160:53]
  wire [31:0] _GEN_23 = _T_235 ? _GEN_18 : 32'h0; // @[ID.scala 160:53]
  wire  _GEN_24 = _T_235 & _GEN_19; // @[ID.scala 160:53]
  wire [31:0] _GEN_25 = _T_235 ? excep_pc : rs1Val; // @[ID.scala 160:53]
  wire [31:0] _GEN_26 = _T_235 ? 32'h4 : _T_234; // @[ID.scala 160:53]
  wire [4:0] _GEN_27 = _T_235 ? 5'h0 : decRes_1; // @[ID.scala 160:53]
  wire  _T_252 = rs1Val < rs2Val; // @[ID.scala 175:35]
  wire [31:0] _T_253 = _T_188 ? 32'h0 : _T_192; // @[ID.scala 175:52]
  wire [31:0] _T_254 = _T_193 ? 32'h0 : _T_197; // @[ID.scala 175:68]
  wire  _T_255 = $signed(_T_253) < $signed(_T_254); // @[ID.scala 175:59]
  wire  _T_256 = decRes_1[0] ? _T_252 : _T_255; // @[ID.scala 175:20]
  wire  _T_258 = rs1Val > rs2Val; // @[ID.scala 176:35]
  wire  _T_261 = $signed(_T_253) > $signed(_T_254); // @[ID.scala 176:59]
  wire  _T_262 = decRes_1[0] ? _T_258 : _T_261; // @[ID.scala 176:20]
  wire  _T_263 = rs1Val == rs2Val; // @[ID.scala 177:24]
  wire  _T_265 = _T_256 & decRes_1[3]; // @[ID.scala 178:23]
  wire  _T_267 = _T_263 & decRes_1[2]; // @[ID.scala 178:37]
  wire  _T_268 = _T_265 | _T_267; // @[ID.scala 178:32]
  wire  _T_270 = _T_262 & decRes_1[1]; // @[ID.scala 178:51]
  wire  _T_271 = _T_268 | _T_270; // @[ID.scala 178:46]
  wire [31:0] _T_283 = excep_pc + _T_234; // @[ID.scala 182:27]
  wire  _T_285 = |_T_283[1:0]; // @[ID.scala 127:22]
  wire [31:0] _GEN_29 = _T_243 ? _T_283 : excep_value; // @[ID.scala 128:26]
  wire  _GEN_31 = _T_285 ? _GEN_12 : excep_valid; // @[ID.scala 127:27]
  wire [31:0] _GEN_32 = _T_285 ? _GEN_29 : excep_value; // @[ID.scala 127:27]
  wire [31:0] _GEN_33 = _T_285 ? _GEN_14 : excep_code; // @[ID.scala 127:27]
  wire [31:0] _GEN_34 = _T_285 ? 32'h0 : _T_283; // @[ID.scala 127:27]
  wire  _GEN_35 = _T_285 ? 1'h0 : 1'h1; // @[ID.scala 127:27]
  wire  _GEN_36 = _T_271 ? _GEN_31 : excep_valid; // @[ID.scala 181:20]
  wire [31:0] _GEN_37 = _T_271 ? _GEN_32 : excep_value; // @[ID.scala 181:20]
  wire [31:0] _GEN_38 = _T_271 ? _GEN_33 : excep_code; // @[ID.scala 181:20]
  wire [31:0] _GEN_39 = _T_271 ? _GEN_34 : 32'h0; // @[ID.scala 181:20]
  wire  _GEN_40 = _T_271 & _GEN_35; // @[ID.scala 181:20]
  wire [31:0] _T_292 = decRes_1[0] ? excep_pc : 32'h0; // @[ID.scala 192:31]
  wire  _T_309 = 4'h7 == decRes_0; // @[Conditional.scala 37:30]
  wire  _T_311 = |inst[14:12]; // @[ID.scala 207:19]
  wire [31:0] _T_314 = inst[14] ? {{27'd0}, rs1Addr} : rs1Val; // @[ID.scala 209:26]
  wire [31:0] _T_315 = csrVal | _T_314; // @[ID.scala 212:33]
  wire [31:0] _T_316 = ~_T_314; // @[ID.scala 213:35]
  wire [31:0] _T_317 = csrVal & _T_316; // @[ID.scala 213:33]
  wire  _T_318 = 2'h1 == inst[13:12]; // @[Mux.scala 80:60]
  wire [31:0] _T_319 = _T_318 ? _T_314 : 32'h0; // @[Mux.scala 80:57]
  wire  _T_320 = 2'h2 == inst[13:12]; // @[Mux.scala 80:60]
  wire [31:0] _T_321 = _T_320 ? _T_315 : _T_319; // @[Mux.scala 80:57]
  wire  _T_322 = 2'h3 == inst[13:12]; // @[Mux.scala 80:60]
  wire [31:0] _T_323 = _T_322 ? _T_317 : _T_321; // @[Mux.scala 80:57]
  wire  _T_325 = inst[31:25] == 7'h9; // @[ID.scala 221:31]
  wire  _T_327 = io_csr_prv >= 2'h1; // @[ID.scala 225:48]
  wire [4:0] _T_329 = _T_188 ? 5'h15 : 5'h14; // @[ID.scala 226:18]
  wire [4:0] _T_330 = _T_327 ? _T_329 : 5'h2; // @[ID.scala 225:36]
  wire [31:0] _GEN_50 = _T_243 ? rs1Val : excep_value; // @[ID.scala 222:30]
  wire [31:0] _GEN_51 = _T_243 ? {{27'd0}, _T_330} : excep_code; // @[ID.scala 222:30]
  wire  _T_333 = 5'h0 == rs2Addr; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_213 = {{2'd0}, io_csr_prv}; // @[Const.scala 131:31]
  wire [3:0] _T_335 = 4'h8 | _GEN_213; // @[Const.scala 131:31]
  wire  _T_336 = 5'h1 == rs2Addr; // @[Conditional.scala 37:30]
  wire  _T_337 = 5'h2 == rs2Addr; // @[Conditional.scala 37:30]
  wire  _T_339 = io_csr_prv >= inst[29:28]; // @[ID.scala 245:52]
  wire [4:0] _GEN_214 = {{3'd0}, inst[29:28]}; // @[Const.scala 132:30]
  wire [4:0] _T_341 = 5'h10 | _GEN_214; // @[Const.scala 132:30]
  wire [4:0] _T_342 = _T_339 ? _T_341 : 5'h2; // @[ID.scala 245:40]
  wire  _GEN_52 = _T_337 | excep_valid; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_53 = _T_337 ? {{27'd0}, _T_342} : excep_code; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_336 | _GEN_52; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_55 = _T_336 ? 32'h3 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_333 | _GEN_54; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_57 = _T_333 ? {{28'd0}, _T_335} : _GEN_55; // @[Conditional.scala 40:58]
  wire  _GEN_58 = _T_243 ? _GEN_56 : excep_valid; // @[ID.scala 232:30]
  wire [31:0] _GEN_59 = _T_243 ? _GEN_57 : excep_code; // @[ID.scala 232:30]
  wire  _GEN_60 = _T_325 ? _GEN_12 : _GEN_58; // @[ID.scala 221:59]
  wire [31:0] _GEN_61 = _T_325 ? _GEN_50 : excep_value; // @[ID.scala 221:59]
  wire [31:0] _GEN_62 = _T_325 ? _GEN_51 : _GEN_59; // @[ID.scala 221:59]
  wire [11:0] _GEN_64 = _T_311 ? csrAddr : 12'h0; // @[ID.scala 207:24]
  wire [31:0] _GEN_65 = _T_311 ? _T_323 : 32'h0; // @[ID.scala 207:24]
  wire [4:0] _GEN_66 = _T_311 ? rdAddr : 5'h0; // @[ID.scala 207:24]
  wire [31:0] _GEN_67 = _T_311 ? csrVal : 32'h0; // @[ID.scala 207:24]
  wire  _GEN_68 = _T_311 ? excep_valid : _GEN_60; // @[ID.scala 207:24]
  wire [31:0] _GEN_69 = _T_311 ? excep_value : _GEN_61; // @[ID.scala 207:24]
  wire [31:0] _GEN_70 = _T_311 ? excep_code : _GEN_62; // @[ID.scala 207:24]
  wire  _T_343 = 4'h8 == decRes_0; // @[Conditional.scala 37:30]
  wire  _T_345 = inst[14:12] == 3'h1; // @[ID.scala 254:26]
  wire  _T_346 = fenceICnt == 2'h3; // @[ID.scala 255:26]
  wire [1:0] _T_348 = fenceICnt + 2'h1; // @[ID.scala 259:36]
  wire  _GEN_72 = _T_346 ? 1'h0 : 1'h1; // @[ID.scala 255:35]
  wire [31:0] _GEN_73 = _T_346 ? 32'h0 : excep_pc; // @[ID.scala 255:35]
  wire  _GEN_75 = _T_345 & _GEN_72; // @[ID.scala 254:40]
  wire [31:0] _GEN_76 = _T_345 ? _GEN_73 : 32'h0; // @[ID.scala 254:40]
  wire  _T_349 = 4'h0 == decRes_0; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_78 = _T_243 ? inst : excep_value; // @[ID.scala 267:28]
  wire [31:0] _GEN_79 = _T_243 ? 32'h2 : excep_code; // @[ID.scala 267:28]
  wire  _GEN_80 = _T_349 ? _GEN_12 : excep_valid; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_81 = _T_349 ? _GEN_78 : excep_value; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_82 = _T_349 ? _GEN_79 : excep_code; // @[Conditional.scala 39:67]
  wire  _GEN_84 = _T_343 & _GEN_75; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_85 = _T_343 ? _GEN_76 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_86 = _T_343 ? excep_valid : _GEN_80; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_87 = _T_343 ? excep_value : _GEN_81; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_88 = _T_343 ? excep_code : _GEN_82; // @[Conditional.scala 39:67]
  wire  _GEN_89 = _T_309 & _T_311; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_90 = _T_309 ? _GEN_64 : 12'h0; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_91 = _T_309 ? _GEN_65 : 32'h0; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_92 = _T_309 ? _GEN_66 : 5'h0; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_93 = _T_309 ? _GEN_67 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_94 = _T_309 ? _GEN_68 : _GEN_86; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_95 = _T_309 ? _GEN_69 : _GEN_87; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_96 = _T_309 ? _GEN_70 : _GEN_88; // @[Conditional.scala 39:67]
  wire  _GEN_98 = _T_309 ? 1'h0 : _GEN_84; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_99 = _T_309 ? 32'h0 : _GEN_85; // @[Conditional.scala 39:67]
  wire  _GEN_101 = _T_293 ? _GEN_31 : _GEN_94; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_102 = _T_293 ? _GEN_32 : _GEN_95; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_103 = _T_293 ? _GEN_33 : _GEN_96; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_104 = _T_293 ? _GEN_34 : _GEN_99; // @[Conditional.scala 39:67]
  wire  _GEN_105 = _T_293 ? _GEN_35 : _GEN_98; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_106 = _T_293 ? excep_pc : _GEN_93; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_107 = _T_293 ? 32'h4 : 32'h0; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_108 = _T_293 ? 5'h0 : decRes_1; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_109 = _T_293 ? rdAddr : _GEN_92; // @[Conditional.scala 39:67]
  wire  _GEN_110 = _T_293 ? 1'h0 : _GEN_89; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_111 = _T_293 ? 12'h0 : _GEN_90; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_112 = _T_293 ? 32'h0 : _GEN_91; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_115 = _T_287 ? _T_234 : _GEN_106; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_116 = _T_287 ? _T_292 : _GEN_107; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_117 = _T_287 ? 5'h0 : _GEN_108; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_118 = _T_287 ? rdAddr : _GEN_109; // @[Conditional.scala 39:67]
  wire  _GEN_119 = _T_287 ? excep_valid : _GEN_101; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_120 = _T_287 ? excep_value : _GEN_102; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_121 = _T_287 ? excep_code : _GEN_103; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_122 = _T_287 ? 32'h0 : _GEN_104; // @[Conditional.scala 39:67]
  wire  _GEN_123 = _T_287 ? 1'h0 : _GEN_105; // @[Conditional.scala 39:67]
  wire  _GEN_124 = _T_287 ? 1'h0 : _GEN_110; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_125 = _T_287 ? 12'h0 : _GEN_111; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_126 = _T_287 ? 32'h0 : _GEN_112; // @[Conditional.scala 39:67]
  wire  _GEN_129 = _T_213 ? _GEN_36 : _GEN_119; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_130 = _T_213 ? _GEN_37 : _GEN_120; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_131 = _T_213 ? _GEN_38 : _GEN_121; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_132 = _T_213 ? _GEN_39 : _GEN_122; // @[Conditional.scala 39:67]
  wire  _GEN_133 = _T_213 ? _GEN_40 : _GEN_123; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_136 = _T_213 ? 32'h0 : _GEN_115; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_137 = _T_213 ? 32'h0 : _GEN_116; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_138 = _T_213 ? decRes_1 : _GEN_117; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_139 = _T_213 ? 5'h0 : _GEN_118; // @[Conditional.scala 39:67]
  wire  _GEN_140 = _T_213 ? 1'h0 : _GEN_124; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_141 = _T_213 ? 12'h0 : _GEN_125; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_142 = _T_213 ? 32'h0 : _GEN_126; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_145 = _T_212 ? rs1Val : _GEN_136; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_146 = _T_212 ? _T_234 : _GEN_137; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_147 = _T_212 ? rs2Val : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_148 = _T_212 ? excep_valid : _GEN_129; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_149 = _T_212 ? excep_value : _GEN_130; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_150 = _T_212 ? excep_code : _GEN_131; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_151 = _T_212 ? 32'h0 : _GEN_132; // @[Conditional.scala 39:67]
  wire  _GEN_152 = _T_212 ? 1'h0 : _GEN_133; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_155 = _T_212 ? decRes_1 : _GEN_138; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_156 = _T_212 ? 5'h0 : _GEN_139; // @[Conditional.scala 39:67]
  wire  _GEN_157 = _T_212 ? 1'h0 : _GEN_140; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_158 = _T_212 ? 12'h0 : _GEN_141; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_159 = _T_212 ? 32'h0 : _GEN_142; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_162 = _T_211 ? _GEN_25 : _GEN_145; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_163 = _T_211 ? _GEN_26 : _GEN_146; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_164 = _T_211 ? rdAddr : _GEN_156; // @[Conditional.scala 39:67]
  wire  _GEN_165 = _T_211 ? _GEN_20 : _GEN_148; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_166 = _T_211 ? _GEN_21 : _GEN_149; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_167 = _T_211 ? _GEN_22 : _GEN_150; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_168 = _T_211 ? _GEN_23 : _GEN_151; // @[Conditional.scala 39:67]
  wire  _GEN_169 = _T_211 ? _GEN_24 : _GEN_152; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_170 = _T_211 ? _GEN_27 : _GEN_155; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_171 = _T_211 ? 32'h0 : _GEN_147; // @[Conditional.scala 39:67]
  wire  _GEN_174 = _T_211 ? 1'h0 : _GEN_157; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_175 = _T_211 ? 12'h0 : _GEN_158; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_176 = _T_211 ? 32'h0 : _GEN_159; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_178 = _T_210 ? rs1Val : _GEN_162; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_179 = _T_210 ? rs2Val : _GEN_163; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_180 = _T_210 ? rdAddr : _GEN_164; // @[Conditional.scala 40:58]
  wire  _GEN_182 = _T_210 ? excep_valid : _GEN_165; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_183 = _T_210 ? excep_value : _GEN_166; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_184 = _T_210 ? excep_code : _GEN_167; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_185 = _T_210 ? 32'h0 : _GEN_168; // @[Conditional.scala 40:58]
  wire  _GEN_186 = _T_210 ? 1'h0 : _GEN_169; // @[Conditional.scala 40:58]
  wire [4:0] _GEN_187 = _T_210 ? decRes_1 : _GEN_170; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_188 = _T_210 ? 32'h0 : _GEN_171; // @[Conditional.scala 40:58]
  wire  _GEN_191 = _T_210 ? 1'h0 : _GEN_174; // @[Conditional.scala 40:58]
  wire [11:0] _GEN_192 = _T_210 ? 12'h0 : _GEN_175; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_193 = _T_210 ? 32'h0 : _GEN_176; // @[Conditional.scala 40:58]
  assign io_iff_branch_valid = stall ? 1'h0 : _GEN_186; // @[ID.scala 102:17 ID.scala 143:25 ID.scala 135:27 ID.scala 135:27 ID.scala 135:27 ID.scala 260:33]
  assign io_iff_branch_bits = stall ? 32'h0 : _GEN_185; // @[ID.scala 102:17 ID.scala 134:26 ID.scala 134:26 ID.scala 134:26 ID.scala 261:32]
  assign io_iff_ready = stall ? 1'h0 : 1'h1; // @[ID.scala 144:18 ID.scala 146:18]
  assign io_reg_read1_addr = inst[19:15]; // @[ID.scala 72:21]
  assign io_reg_read2_addr = inst[24:20]; // @[ID.scala 73:21]
  assign io_ex_aluOp_rd1 = stall ? 32'h0 : _GEN_178; // @[ID.scala 103:15 ID.scala 150:25 ID.scala 156:25 ID.scala 162:27 ID.scala 169:25 ID.scala 190:25 ID.scala 199:25 ID.scala 219:30]
  assign io_ex_aluOp_rd2 = stall ? 32'h0 : _GEN_179; // @[ID.scala 103:15 ID.scala 151:25 ID.scala 157:25 ID.scala 163:27 ID.scala 170:25 ID.scala 192:25 ID.scala 200:25]
  assign io_ex_aluOp_opt = stall ? 5'h0 : _GEN_187; // @[ID.scala 103:15 ID.scala 104:19 ID.scala 142:21 ID.scala 164:27 ID.scala 193:27 ID.scala 201:25]
  assign io_ex_wrRegOp_addr = stall ? 5'h0 : _GEN_180; // @[ID.scala 106:17 ID.scala 141:24 ID.scala 152:28 ID.scala 158:28 ID.scala 194:28 ID.scala 202:28 ID.scala 218:30]
  assign io_ex_wrCSROp_valid = stall ? 1'h0 : _GEN_191; // @[ID.scala 105:17 ID.scala 215:31]
  assign io_ex_wrCSROp_addr = stall ? 12'h0 : _GEN_192; // @[ID.scala 105:17 ID.scala 216:30]
  assign io_ex_wrCSROp_data = stall ? 32'h0 : _GEN_193; // @[ID.scala 105:17 ID.scala 217:30]
  assign io_ex_store_data = stall ? 32'h0 : _GEN_188; // @[ID.scala 109:20 ID.scala 171:26]
  assign io_ex_excep_valid = stall ? excep_valid : _GEN_182; // @[ID.scala 107:15 ID.scala 129:27 ID.scala 129:27 ID.scala 129:27 ID.scala 223:31 ID.scala 235:35 ID.scala 239:35 ID.scala 244:35 ID.scala 268:29]
  assign io_ex_excep_code = stall ? excep_code : _GEN_184; // @[ID.scala 107:15 ID.scala 131:26 ID.scala 131:26 ID.scala 131:26 ID.scala 225:30 ID.scala 236:34 ID.scala 240:34 ID.scala 245:34 ID.scala 270:28]
  assign io_ex_excep_value = stall ? excep_value : _GEN_183; // @[ID.scala 107:15 ID.scala 130:27 ID.scala 130:27 ID.scala 130:27 ID.scala 224:31 ID.scala 269:29]
  assign io_ex_excep_pc = excep_pc; // @[ID.scala 107:15]
  assign io_ex_excep_valid_inst = excep_valid_inst & _T_207; // @[ID.scala 107:15 ID.scala 108:26]
  assign io_csr_addr = inst[31:20]; // @[ID.scala 74:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  excep_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  excep_code = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  excep_value = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  excep_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  excep_valid_inst = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  fenceICnt = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      inst <= 32'h13;
    end else if (io_flush) begin
      inst <= 32'h13;
    end else if (!(stall)) begin
      inst <= io_iff_inst;
    end
    if (reset) begin
      excep_valid <= 1'h0;
    end else if (io_flush) begin
      excep_valid <= 1'h0;
    end else if (!(stall)) begin
      excep_valid <= io_iff_excep_valid;
    end
    if (reset) begin
      excep_code <= 32'h0;
    end else if (io_flush) begin
      excep_code <= 32'h0;
    end else if (!(stall)) begin
      excep_code <= io_iff_excep_code;
    end
    if (reset) begin
      excep_value <= 32'h0;
    end else if (io_flush) begin
      excep_value <= 32'h0;
    end else if (!(stall)) begin
      excep_value <= io_iff_excep_value;
    end
    if (reset) begin
      excep_pc <= 32'h0;
    end else if (io_flush) begin
      excep_pc <= 32'h0;
    end else if (!(stall)) begin
      excep_pc <= io_iff_excep_pc;
    end
    if (reset) begin
      excep_valid_inst <= 1'h0;
    end else if (io_flush) begin
      excep_valid_inst <= 1'h0;
    end else if (!(stall)) begin
      excep_valid_inst <= io_iff_excep_valid_inst;
    end
    if (reset) begin
      fenceICnt <= 2'h0;
    end else if (!(stall)) begin
      if (!(_T_210)) begin
        if (!(_T_211)) begin
          if (!(_T_212)) begin
            if (!(_T_213)) begin
              if (!(_T_287)) begin
                if (!(_T_293)) begin
                  if (!(_T_309)) begin
                    if (_T_343) begin
                      if (_T_345) begin
                        if (_T_346) begin
                          fenceICnt <= 2'h0;
                        end else begin
                          fenceICnt <= _T_348;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module EX(
  input         clock,
  input         reset,
  input  [31:0] io_id_aluOp_rd1,
  input  [31:0] io_id_aluOp_rd2,
  input  [4:0]  io_id_aluOp_opt,
  input  [4:0]  io_id_wrRegOp_addr,
  input         io_id_wrCSROp_valid,
  input  [11:0] io_id_wrCSROp_addr,
  input  [31:0] io_id_wrCSROp_data,
  input  [31:0] io_id_store_data,
  input         io_id_excep_valid,
  input  [31:0] io_id_excep_code,
  input  [31:0] io_id_excep_value,
  input  [31:0] io_id_excep_pc,
  input         io_id_excep_valid_inst,
  output        io_id_ready,
  output [31:0] io_mem_ramOp_addr,
  output [3:0]  io_mem_ramOp_mode,
  output [31:0] io_mem_ramOp_wdata,
  output [4:0]  io_mem_wrRegOp_addr,
  output [31:0] io_mem_wrRegOp_data,
  output        io_mem_wrRegOp_rdy,
  output        io_mem_wrCSROp_valid,
  output [11:0] io_mem_wrCSROp_addr,
  output [31:0] io_mem_wrCSROp_data,
  output        io_mem_excep_valid,
  output [31:0] io_mem_excep_code,
  output [31:0] io_mem_excep_value,
  output [31:0] io_mem_excep_pc,
  output        io_mem_excep_valid_inst,
  input         io_mem_ready,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] alu_rd1; // @[EX.scala 18:20]
  reg [31:0] alu_rd2; // @[EX.scala 18:20]
  reg [4:0] alu_opt; // @[EX.scala 18:20]
  wire [4:0] shamt = alu_rd2[4:0]; // @[EX.scala 24:16]
  wire [31:0] _T_2 = alu_rd1 + alu_rd2; // @[EX.scala 28:7]
  wire [31:0] _T_6 = alu_rd1 - alu_rd2; // @[EX.scala 31:17]
  wire [31:0] _T_7 = alu_rd1; // @[EX.scala 32:20]
  wire  _T_9 = $signed(alu_rd1) < $signed(alu_rd2); // @[EX.scala 32:27]
  wire  _T_11 = alu_rd1 < alu_rd2; // @[EX.scala 33:21]
  wire [31:0] _T_13 = alu_rd1 ^ alu_rd2; // @[EX.scala 34:17]
  wire [31:0] _T_14 = alu_rd1 | alu_rd2; // @[EX.scala 35:16]
  wire [31:0] _T_15 = alu_rd1 & alu_rd2; // @[EX.scala 36:17]
  wire [62:0] _GEN_20 = {{31'd0}, alu_rd1}; // @[EX.scala 37:17]
  wire [62:0] _T_16 = _GEN_20 << shamt; // @[EX.scala 37:17]
  wire [31:0] _T_17 = alu_rd1 >> shamt; // @[EX.scala 38:17]
  wire [31:0] _T_20 = $signed(alu_rd1) >>> shamt; // @[EX.scala 39:34]
  wire [63:0] _T_21 = alu_rd1 * alu_rd2; // @[EX.scala 41:17]
  wire [63:0] _T_25 = $signed(alu_rd1) * $signed(alu_rd2); // @[EX.scala 42:25]
  wire [32:0] _T_30 = {1'b0,$signed(alu_rd2)}; // @[EX.scala 44:27]
  wire [32:0] _GEN_21 = {{1{_T_7[31]}},_T_7}; // @[EX.scala 44:27]
  wire [64:0] _T_31 = $signed(_GEN_21) * $signed(_T_30); // @[EX.scala 44:27]
  wire [63:0] _T_33 = _T_31[63:0]; // @[EX.scala 44:27]
  wire [32:0] _T_38 = $signed(alu_rd1) / $signed(alu_rd2); // @[EX.scala 45:36]
  wire [31:0] _T_39 = alu_rd1 / alu_rd2; // @[EX.scala 46:17]
  wire [31:0] _T_43 = $signed(alu_rd1) % $signed(alu_rd2); // @[EX.scala 47:37]
  wire [31:0] _GEN_0 = alu_rd1 % alu_rd2; // @[EX.scala 48:17]
  wire [31:0] _T_44 = _GEN_0[31:0]; // @[EX.scala 48:17]
  wire  _T_45 = 5'h0 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_46 = _T_45 ? _T_2 : _T_2; // @[Mux.scala 80:57]
  wire  _T_47 = 5'h1 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_48 = _T_47 ? _T_6 : _T_46; // @[Mux.scala 80:57]
  wire  _T_49 = 5'h2 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_50 = _T_49 ? {{31'd0}, _T_9} : _T_48; // @[Mux.scala 80:57]
  wire  _T_51 = 5'h3 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_52 = _T_51 ? {{31'd0}, _T_11} : _T_50; // @[Mux.scala 80:57]
  wire  _T_53 = 5'h4 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_54 = _T_53 ? _T_13 : _T_52; // @[Mux.scala 80:57]
  wire  _T_55 = 5'h5 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_56 = _T_55 ? _T_14 : _T_54; // @[Mux.scala 80:57]
  wire  _T_57 = 5'h6 == alu_opt; // @[Mux.scala 80:60]
  wire [31:0] _T_58 = _T_57 ? _T_15 : _T_56; // @[Mux.scala 80:57]
  wire  _T_59 = 5'h7 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_60 = _T_59 ? _T_16 : {{31'd0}, _T_58}; // @[Mux.scala 80:57]
  wire  _T_61 = 5'h8 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_62 = _T_61 ? {{31'd0}, _T_17} : _T_60; // @[Mux.scala 80:57]
  wire  _T_63 = 5'h9 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_64 = _T_63 ? {{31'd0}, _T_20} : _T_62; // @[Mux.scala 80:57]
  wire  _T_65 = 5'hb == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_66 = _T_65 ? {{31'd0}, _T_21[31:0]} : _T_64; // @[Mux.scala 80:57]
  wire  _T_67 = 5'hc == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_68 = _T_67 ? {{31'd0}, _T_25[63:32]} : _T_66; // @[Mux.scala 80:57]
  wire  _T_69 = 5'he == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_70 = _T_69 ? {{31'd0}, _T_21[63:32]} : _T_68; // @[Mux.scala 80:57]
  wire  _T_71 = 5'hd == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_72 = _T_71 ? {{31'd0}, _T_33[63:32]} : _T_70; // @[Mux.scala 80:57]
  wire  _T_73 = 5'hf == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_74 = _T_73 ? {{30'd0}, _T_38} : _T_72; // @[Mux.scala 80:57]
  wire  _T_75 = 5'h10 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_76 = _T_75 ? {{31'd0}, _T_39} : _T_74; // @[Mux.scala 80:57]
  wire  _T_77 = 5'h11 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] _T_78 = _T_77 ? {{31'd0}, _T_43} : _T_76; // @[Mux.scala 80:57]
  wire  _T_79 = 5'h12 == alu_opt; // @[Mux.scala 80:60]
  wire [62:0] aluRes = _T_79 ? {{31'd0}, _T_44} : _T_78; // @[Mux.scala 80:57]
  reg [4:0] wregAddr; // @[EX.scala 56:27]
  reg [31:0] store_data; // @[EX.scala 57:27]
  wire [4:0] _T_80 = alu_opt & 5'h18; // @[EX.scala 61:31]
  wire  _T_82 = 5'h18 == alu_opt; // @[Mux.scala 80:60]
  wire  _T_84 = 5'h1c == alu_opt; // @[Mux.scala 80:60]
  wire [2:0] _T_85 = _T_84 ? 3'h4 : {{2'd0}, _T_82}; // @[Mux.scala 80:57]
  wire  _T_86 = 5'h1d == alu_opt; // @[Mux.scala 80:60]
  wire [2:0] _T_87 = _T_86 ? 3'h5 : _T_85; // @[Mux.scala 80:57]
  wire  _T_88 = 5'h1a == alu_opt; // @[Mux.scala 80:60]
  wire [2:0] _T_89 = _T_88 ? 3'h2 : _T_87; // @[Mux.scala 80:57]
  wire  _T_90 = 5'h1b == alu_opt; // @[Mux.scala 80:60]
  wire [2:0] _T_91 = _T_90 ? 3'h3 : _T_89; // @[Mux.scala 80:57]
  wire  _T_92 = 5'h14 == alu_opt; // @[Mux.scala 80:60]
  wire [3:0] _T_93 = _T_92 ? 4'h9 : {{1'd0}, _T_91}; // @[Mux.scala 80:57]
  wire  _T_94 = 5'h15 == alu_opt; // @[Mux.scala 80:60]
  wire [3:0] _T_95 = _T_94 ? 4'ha : _T_93; // @[Mux.scala 80:57]
  wire  _T_96 = 5'h16 == alu_opt; // @[Mux.scala 80:60]
  reg  excep_valid; // @[EX.scala 78:24]
  reg [31:0] excep_code; // @[EX.scala 78:24]
  reg [31:0] excep_value; // @[EX.scala 78:24]
  reg [31:0] excep_pc; // @[EX.scala 78:24]
  reg  excep_valid_inst; // @[EX.scala 78:24]
  reg  wrCSROp_valid; // @[EX.scala 79:24]
  reg [11:0] wrCSROp_addr; // @[EX.scala 79:24]
  reg [31:0] wrCSROp_data; // @[EX.scala 79:24]
  reg [2:0] countdown; // @[EX.scala 85:26]
  wire  _T_98 = ~io_mem_ready; // @[EX.scala 87:15]
  wire  _T_99 = countdown != 3'h0; // @[EX.scala 87:42]
  wire  stall = _T_98 | _T_99; // @[EX.scala 87:29]
  wire  _T_100 = ~stall; // @[EX.scala 89:18]
  wire  _T_102 = io_id_aluOp_opt >= 5'hb; // @[EX.scala 92:34]
  wire  _T_103 = _T_100 & _T_102; // @[EX.scala 92:15]
  wire  _T_104 = io_id_aluOp_opt <= 5'h12; // @[EX.scala 92:61]
  wire  _T_105 = _T_103 & _T_104; // @[EX.scala 92:42]
  wire [2:0] _T_108 = countdown - 3'h1; // @[EX.scala 95:28]
  assign io_id_ready = ~stall; // @[EX.scala 89:15]
  assign io_mem_ramOp_addr = aluRes[31:0]; // @[EX.scala 63:21]
  assign io_mem_ramOp_mode = _T_96 ? 4'hc : _T_95; // @[EX.scala 64:21]
  assign io_mem_ramOp_wdata = store_data; // @[EX.scala 74:22]
  assign io_mem_wrRegOp_addr = wregAddr; // @[EX.scala 59:23]
  assign io_mem_wrRegOp_data = aluRes[31:0]; // @[EX.scala 60:23]
  assign io_mem_wrRegOp_rdy = _T_80 != 5'h18; // @[EX.scala 61:23]
  assign io_mem_wrCSROp_valid = wrCSROp_valid; // @[EX.scala 81:18]
  assign io_mem_wrCSROp_addr = wrCSROp_addr; // @[EX.scala 81:18]
  assign io_mem_wrCSROp_data = wrCSROp_data; // @[EX.scala 81:18]
  assign io_mem_excep_valid = excep_valid; // @[EX.scala 80:18]
  assign io_mem_excep_code = excep_code; // @[EX.scala 80:18]
  assign io_mem_excep_value = excep_value; // @[EX.scala 80:18]
  assign io_mem_excep_pc = excep_pc; // @[EX.scala 80:18]
  assign io_mem_excep_valid_inst = excep_valid_inst; // @[EX.scala 80:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alu_rd1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  alu_rd2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  alu_opt = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  wregAddr = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  store_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  excep_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  excep_code = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  excep_value = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  excep_pc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  excep_valid_inst = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  wrCSROp_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  wrCSROp_addr = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  wrCSROp_data = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  countdown = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      alu_rd1 <= 32'h0;
    end else if (!(stall)) begin
      alu_rd1 <= io_id_aluOp_rd1;
    end
    if (reset) begin
      alu_rd2 <= 32'h0;
    end else if (!(stall)) begin
      alu_rd2 <= io_id_aluOp_rd2;
    end
    if (reset) begin
      alu_opt <= 5'h0;
    end else if (io_flush) begin
      alu_opt <= 5'h0;
    end else if (!(stall)) begin
      alu_opt <= io_id_aluOp_opt;
    end
    if (reset) begin
      wregAddr <= 5'h0;
    end else if (io_flush) begin
      wregAddr <= 5'h0;
    end else if (!(stall)) begin
      wregAddr <= io_id_wrRegOp_addr;
    end
    if (reset) begin
      store_data <= 32'h0;
    end else if (!(stall)) begin
      store_data <= io_id_store_data;
    end
    if (io_flush) begin
      excep_valid <= 1'h0;
    end else if (!(stall)) begin
      excep_valid <= io_id_excep_valid;
    end
    if (!(stall)) begin
      excep_code <= io_id_excep_code;
    end
    if (!(stall)) begin
      excep_value <= io_id_excep_value;
    end
    if (!(stall)) begin
      excep_pc <= io_id_excep_pc;
    end
    if (io_flush) begin
      excep_valid_inst <= 1'h0;
    end else if (!(stall)) begin
      excep_valid_inst <= io_id_excep_valid_inst;
    end
    if (io_flush) begin
      wrCSROp_valid <= 1'h0;
    end else if (!(stall)) begin
      wrCSROp_valid <= io_id_wrCSROp_valid;
    end
    if (!(stall)) begin
      wrCSROp_addr <= io_id_wrCSROp_addr;
    end
    if (!(stall)) begin
      wrCSROp_data <= io_id_wrCSROp_data;
    end
    if (reset) begin
      countdown <= 3'h0;
    end else if (_T_105) begin
      countdown <= 3'h7;
    end else if (_T_99) begin
      countdown <= _T_108;
    end else begin
      countdown <= 3'h0;
    end
  end
endmodule
module MEM(
  input         clock,
  input         reset,
  input  [31:0] io_ex_ramOp_addr,
  input  [3:0]  io_ex_ramOp_mode,
  input  [31:0] io_ex_ramOp_wdata,
  input  [4:0]  io_ex_wrRegOp_addr,
  input  [31:0] io_ex_wrRegOp_data,
  input         io_ex_wrCSROp_valid,
  input  [11:0] io_ex_wrCSROp_addr,
  input  [31:0] io_ex_wrCSROp_data,
  input         io_ex_excep_valid,
  input  [31:0] io_ex_excep_code,
  input  [31:0] io_ex_excep_value,
  input  [31:0] io_ex_excep_pc,
  input         io_ex_excep_valid_inst,
  output        io_ex_ready,
  output [31:0] io_mmu_addr,
  output [3:0]  io_mmu_mode,
  output [31:0] io_mmu_wdata,
  input  [31:0] io_mmu_rdata,
  input         io_mmu_ok,
  input         io_mmu_pageFault,
  output        io_csr_wrCSROp_valid,
  output [11:0] io_csr_wrCSROp_addr,
  output [31:0] io_csr_wrCSROp_data,
  output        io_csr_excep_valid,
  output [31:0] io_csr_excep_code,
  output [31:0] io_csr_excep_value,
  output [31:0] io_csr_excep_pc,
  output        io_csr_excep_valid_inst,
  input         io_csr_inter_valid,
  input  [31:0] io_csr_inter_bits,
  output [4:0]  io_reg_addr,
  output [31:0] io_reg_data,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ramOp_addr; // @[MEM.scala 17:24]
  reg [3:0] ramOp_mode; // @[MEM.scala 17:24]
  reg [31:0] ramOp_wdata; // @[MEM.scala 17:24]
  reg [4:0] reg_addr; // @[MEM.scala 18:24]
  reg [31:0] reg_data; // @[MEM.scala 18:24]
  reg  wrCSROp_valid; // @[MEM.scala 19:24]
  reg [11:0] wrCSROp_addr; // @[MEM.scala 19:24]
  reg [31:0] wrCSROp_data; // @[MEM.scala 19:24]
  reg  excep_valid; // @[MEM.scala 20:24]
  reg [31:0] excep_code; // @[MEM.scala 20:24]
  reg [31:0] excep_value; // @[MEM.scala 20:24]
  reg [31:0] excep_pc; // @[MEM.scala 20:24]
  reg  excep_valid_inst; // @[MEM.scala 20:24]
  wire  _T_4 = io_mmu_mode != 4'h0; // @[MEM.scala 23:27]
  wire  _T_5 = ~io_mmu_ok; // @[MEM.scala 23:46]
  wire  stall = _T_4 & _T_5; // @[MEM.scala 23:43]
  wire  _T_6 = ~stall; // @[MEM.scala 24:18]
  wire  _T_8 = io_csr_inter_valid & io_ex_excep_valid_inst; // @[MEM.scala 32:29]
  wire  _GEN_0 = _T_8 | io_ex_excep_valid; // @[MEM.scala 32:56]
  wire  _T_10 = ~ramOp_mode[3]; // @[Const.scala 23:32]
  wire  _T_11 = |ramOp_mode; // @[Const.scala 23:43]
  wire  _T_12 = _T_10 & _T_11; // @[Const.scala 23:38]
  wire  _T_14 = ~excep_valid; // @[MEM.scala 53:8]
  wire  _T_17 = ramOp_mode[1] & ramOp_addr[0]; // @[Bundles.scala 48:24]
  wire  _T_19 = ramOp_mode[2:0] == 3'h1; // @[Const.scala 25:39]
  wire  _T_21 = |ramOp_addr[1:0]; // @[Bundles.scala 49:37]
  wire  _T_22 = _T_19 & _T_21; // @[Bundles.scala 49:24]
  wire  _T_23 = _T_17 | _T_22; // @[Bundles.scala 48:35]
  wire [2:0] _T_28 = _T_12 ? 3'h4 : 3'h6; // @[MEM.scala 60:31]
  wire [3:0] _GEN_16 = _T_23 ? 4'h0 : ramOp_mode; // @[MEM.scala 56:28]
  wire  _GEN_17 = _T_23 | excep_valid; // @[MEM.scala 56:28]
  wire [31:0] _GEN_18 = _T_23 ? ramOp_addr : excep_value; // @[MEM.scala 56:28]
  wire [31:0] _GEN_19 = _T_23 ? {{29'd0}, _T_28} : excep_code; // @[MEM.scala 56:28]
  wire [3:0] _T_33 = _T_12 ? 4'hd : 4'hf; // @[MEM.scala 67:31]
  wire  _GEN_20 = io_mmu_pageFault | _GEN_17; // @[MEM.scala 64:28]
  wire [31:0] _GEN_21 = io_mmu_pageFault ? ramOp_addr : _GEN_18; // @[MEM.scala 64:28]
  wire [31:0] _GEN_22 = io_mmu_pageFault ? {{28'd0}, _T_33} : _GEN_19; // @[MEM.scala 64:28]
  wire [3:0] _GEN_23 = _T_14 ? _GEN_16 : ramOp_mode; // @[MEM.scala 53:22]
  wire  _GEN_24 = _T_14 ? _GEN_20 : excep_valid; // @[MEM.scala 53:22]
  wire [4:0] _GEN_27 = io_csr_excep_valid ? 5'h0 : reg_addr; // @[MEM.scala 74:28]
  wire  _GEN_28 = io_csr_excep_valid ? 1'h0 : wrCSROp_valid; // @[MEM.scala 74:28]
  assign io_ex_ready = ~stall; // @[MEM.scala 24:15]
  assign io_mmu_addr = ramOp_addr; // @[MEM.scala 41:16]
  assign io_mmu_mode = excep_valid ? 4'h0 : _GEN_23; // @[MEM.scala 43:16 MEM.scala 57:19 MEM.scala 81:17]
  assign io_mmu_wdata = ramOp_wdata; // @[MEM.scala 42:16]
  assign io_csr_wrCSROp_valid = stall ? 1'h0 : _GEN_28; // @[MEM.scala 49:18 MEM.scala 76:26 MEM.scala 88:26]
  assign io_csr_wrCSROp_addr = wrCSROp_addr; // @[MEM.scala 49:18]
  assign io_csr_wrCSROp_data = wrCSROp_data; // @[MEM.scala 49:18]
  assign io_csr_excep_valid = stall ? 1'h0 : _GEN_24; // @[MEM.scala 50:16 MEM.scala 58:26 MEM.scala 65:26 MEM.scala 87:24]
  assign io_csr_excep_code = _T_14 ? _GEN_22 : excep_code; // @[MEM.scala 50:16 MEM.scala 60:25 MEM.scala 67:25]
  assign io_csr_excep_value = _T_14 ? _GEN_21 : excep_value; // @[MEM.scala 50:16 MEM.scala 59:26 MEM.scala 66:26]
  assign io_csr_excep_pc = excep_pc; // @[MEM.scala 50:16]
  assign io_csr_excep_valid_inst = stall ? 1'h0 : excep_valid_inst; // @[MEM.scala 50:16 MEM.scala 86:29]
  assign io_reg_addr = stall ? 5'h0 : _GEN_27; // @[MEM.scala 45:15 MEM.scala 75:17 MEM.scala 89:17]
  assign io_reg_data = _T_12 ? io_mmu_rdata : reg_data; // @[MEM.scala 47:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ramOp_addr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ramOp_mode = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  ramOp_wdata = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_addr = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  reg_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  wrCSROp_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  wrCSROp_addr = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  wrCSROp_data = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  excep_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  excep_code = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  excep_value = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  excep_pc = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  excep_valid_inst = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ramOp_addr <= 32'h0;
    end else if (_T_6) begin
      ramOp_addr <= io_ex_ramOp_addr;
    end
    if (reset) begin
      ramOp_mode <= 4'h0;
    end else if (io_flush) begin
      ramOp_mode <= 4'h0;
    end else if (_T_6) begin
      ramOp_mode <= io_ex_ramOp_mode;
    end
    if (reset) begin
      ramOp_wdata <= 32'h0;
    end else if (_T_6) begin
      ramOp_wdata <= io_ex_ramOp_wdata;
    end
    if (reset) begin
      reg_addr <= 5'h0;
    end else if (io_flush) begin
      reg_addr <= 5'h0;
    end else if (_T_6) begin
      reg_addr <= io_ex_wrRegOp_addr;
    end
    if (reset) begin
      reg_data <= 32'h0;
    end else if (_T_6) begin
      reg_data <= io_ex_wrRegOp_data;
    end
    if (reset) begin
      wrCSROp_valid <= 1'h0;
    end else if (io_flush) begin
      wrCSROp_valid <= 1'h0;
    end else if (_T_6) begin
      wrCSROp_valid <= io_ex_wrCSROp_valid;
    end
    if (reset) begin
      wrCSROp_addr <= 12'h0;
    end else if (_T_6) begin
      wrCSROp_addr <= io_ex_wrCSROp_addr;
    end
    if (reset) begin
      wrCSROp_data <= 32'h0;
    end else if (_T_6) begin
      wrCSROp_data <= io_ex_wrCSROp_data;
    end
    if (reset) begin
      excep_valid <= 1'h0;
    end else if (io_flush) begin
      excep_valid <= 1'h0;
    end else if (_T_6) begin
      excep_valid <= _GEN_0;
    end
    if (reset) begin
      excep_code <= 32'h0;
    end else if (_T_6) begin
      if (_T_8) begin
        excep_code <= io_csr_inter_bits;
      end else begin
        excep_code <= io_ex_excep_code;
      end
    end
    if (reset) begin
      excep_value <= 32'h0;
    end else if (_T_6) begin
      excep_value <= io_ex_excep_value;
    end
    if (reset) begin
      excep_pc <= 32'h0;
    end else if (_T_6) begin
      excep_pc <= io_ex_excep_pc;
    end
    if (reset) begin
      excep_valid_inst <= 1'h0;
    end else if (io_flush) begin
      excep_valid_inst <= 1'h0;
    end else if (_T_6) begin
      excep_valid_inst <= io_ex_excep_valid_inst;
    end
  end
endmodule
module RegFile(
  input         clock,
  input  [4:0]  io_id_read1_addr,
  output [31:0] io_id_read1_data,
  input  [4:0]  io_id_read2_addr,
  output [31:0] io_id_read2_data,
  input  [4:0]  io_mem_addr,
  input  [31:0] io_mem_data,
  output [31:0] io_log_0,
  output [31:0] io_log_1,
  output [31:0] io_log_2,
  output [31:0] io_log_3,
  output [31:0] io_log_4,
  output [31:0] io_log_5,
  output [31:0] io_log_6,
  output [31:0] io_log_7,
  output [31:0] io_log_8,
  output [31:0] io_log_9,
  output [31:0] io_log_10,
  output [31:0] io_log_11,
  output [31:0] io_log_12,
  output [31:0] io_log_13,
  output [31:0] io_log_14,
  output [31:0] io_log_15,
  output [31:0] io_log_16,
  output [31:0] io_log_17,
  output [31:0] io_log_18,
  output [31:0] io_log_19,
  output [31:0] io_log_20,
  output [31:0] io_log_21,
  output [31:0] io_log_22,
  output [31:0] io_log_23,
  output [31:0] io_log_24,
  output [31:0] io_log_25,
  output [31:0] io_log_26,
  output [31:0] io_log_27,
  output [31:0] io_log_28,
  output [31:0] io_log_29,
  output [31:0] io_log_30,
  output [31:0] io_log_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] regs [0:31]; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_1_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_1_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_2_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_2_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_5_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_5_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_6_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_6_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_7_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_7_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_8_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_8_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_9_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_9_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_10_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_10_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_11_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_11_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_12_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_12_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_13_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_13_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_14_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_14_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_15_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_15_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_16_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_16_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_17_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_17_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_18_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_18_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_19_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_19_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_20_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_20_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_21_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_21_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_22_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_22_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_23_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_23_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_24_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_24_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_25_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_25_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_26_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_26_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_27_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_27_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_28_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_28_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_29_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_29_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_30_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_30_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_31_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_31_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_32_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_32_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_33_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_33_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_34_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_34_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_35_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_35_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_36_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_36_addr; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_addr; // @[RegFile.scala 14:17]
  wire  regs__T_mask; // @[RegFile.scala 14:17]
  wire  regs__T_en; // @[RegFile.scala 14:17]
  wire [31:0] regs__T_4_data; // @[RegFile.scala 14:17]
  wire [4:0] regs__T_4_addr; // @[RegFile.scala 14:17]
  wire  regs__T_4_mask; // @[RegFile.scala 14:17]
  wire  regs__T_4_en; // @[RegFile.scala 14:17]
  assign regs__T_1_addr = io_id_read1_addr;
  assign regs__T_1_data = regs[regs__T_1_addr]; // @[RegFile.scala 14:17]
  assign regs__T_2_addr = io_id_read2_addr;
  assign regs__T_2_data = regs[regs__T_2_addr]; // @[RegFile.scala 14:17]
  assign regs__T_5_addr = 5'h0;
  assign regs__T_5_data = regs[regs__T_5_addr]; // @[RegFile.scala 14:17]
  assign regs__T_6_addr = 5'h1;
  assign regs__T_6_data = regs[regs__T_6_addr]; // @[RegFile.scala 14:17]
  assign regs__T_7_addr = 5'h2;
  assign regs__T_7_data = regs[regs__T_7_addr]; // @[RegFile.scala 14:17]
  assign regs__T_8_addr = 5'h3;
  assign regs__T_8_data = regs[regs__T_8_addr]; // @[RegFile.scala 14:17]
  assign regs__T_9_addr = 5'h4;
  assign regs__T_9_data = regs[regs__T_9_addr]; // @[RegFile.scala 14:17]
  assign regs__T_10_addr = 5'h5;
  assign regs__T_10_data = regs[regs__T_10_addr]; // @[RegFile.scala 14:17]
  assign regs__T_11_addr = 5'h6;
  assign regs__T_11_data = regs[regs__T_11_addr]; // @[RegFile.scala 14:17]
  assign regs__T_12_addr = 5'h7;
  assign regs__T_12_data = regs[regs__T_12_addr]; // @[RegFile.scala 14:17]
  assign regs__T_13_addr = 5'h8;
  assign regs__T_13_data = regs[regs__T_13_addr]; // @[RegFile.scala 14:17]
  assign regs__T_14_addr = 5'h9;
  assign regs__T_14_data = regs[regs__T_14_addr]; // @[RegFile.scala 14:17]
  assign regs__T_15_addr = 5'ha;
  assign regs__T_15_data = regs[regs__T_15_addr]; // @[RegFile.scala 14:17]
  assign regs__T_16_addr = 5'hb;
  assign regs__T_16_data = regs[regs__T_16_addr]; // @[RegFile.scala 14:17]
  assign regs__T_17_addr = 5'hc;
  assign regs__T_17_data = regs[regs__T_17_addr]; // @[RegFile.scala 14:17]
  assign regs__T_18_addr = 5'hd;
  assign regs__T_18_data = regs[regs__T_18_addr]; // @[RegFile.scala 14:17]
  assign regs__T_19_addr = 5'he;
  assign regs__T_19_data = regs[regs__T_19_addr]; // @[RegFile.scala 14:17]
  assign regs__T_20_addr = 5'hf;
  assign regs__T_20_data = regs[regs__T_20_addr]; // @[RegFile.scala 14:17]
  assign regs__T_21_addr = 5'h10;
  assign regs__T_21_data = regs[regs__T_21_addr]; // @[RegFile.scala 14:17]
  assign regs__T_22_addr = 5'h11;
  assign regs__T_22_data = regs[regs__T_22_addr]; // @[RegFile.scala 14:17]
  assign regs__T_23_addr = 5'h12;
  assign regs__T_23_data = regs[regs__T_23_addr]; // @[RegFile.scala 14:17]
  assign regs__T_24_addr = 5'h13;
  assign regs__T_24_data = regs[regs__T_24_addr]; // @[RegFile.scala 14:17]
  assign regs__T_25_addr = 5'h14;
  assign regs__T_25_data = regs[regs__T_25_addr]; // @[RegFile.scala 14:17]
  assign regs__T_26_addr = 5'h15;
  assign regs__T_26_data = regs[regs__T_26_addr]; // @[RegFile.scala 14:17]
  assign regs__T_27_addr = 5'h16;
  assign regs__T_27_data = regs[regs__T_27_addr]; // @[RegFile.scala 14:17]
  assign regs__T_28_addr = 5'h17;
  assign regs__T_28_data = regs[regs__T_28_addr]; // @[RegFile.scala 14:17]
  assign regs__T_29_addr = 5'h18;
  assign regs__T_29_data = regs[regs__T_29_addr]; // @[RegFile.scala 14:17]
  assign regs__T_30_addr = 5'h19;
  assign regs__T_30_data = regs[regs__T_30_addr]; // @[RegFile.scala 14:17]
  assign regs__T_31_addr = 5'h1a;
  assign regs__T_31_data = regs[regs__T_31_addr]; // @[RegFile.scala 14:17]
  assign regs__T_32_addr = 5'h1b;
  assign regs__T_32_data = regs[regs__T_32_addr]; // @[RegFile.scala 14:17]
  assign regs__T_33_addr = 5'h1c;
  assign regs__T_33_data = regs[regs__T_33_addr]; // @[RegFile.scala 14:17]
  assign regs__T_34_addr = 5'h1d;
  assign regs__T_34_data = regs[regs__T_34_addr]; // @[RegFile.scala 14:17]
  assign regs__T_35_addr = 5'h1e;
  assign regs__T_35_data = regs[regs__T_35_addr]; // @[RegFile.scala 14:17]
  assign regs__T_36_addr = 5'h1f;
  assign regs__T_36_data = regs[regs__T_36_addr]; // @[RegFile.scala 14:17]
  assign regs__T_data = 32'h0;
  assign regs__T_addr = 5'h0;
  assign regs__T_mask = 1'h1;
  assign regs__T_en = 1'h1;
  assign regs__T_4_data = io_mem_data;
  assign regs__T_4_addr = io_mem_addr;
  assign regs__T_4_mask = 1'h1;
  assign regs__T_4_en = |io_mem_addr;
  assign io_id_read1_data = regs__T_1_data; // @[RegFile.scala 20:20]
  assign io_id_read2_data = regs__T_2_data; // @[RegFile.scala 21:20]
  assign io_log_0 = regs__T_5_data; // @[RegFile.scala 32:15]
  assign io_log_1 = regs__T_6_data; // @[RegFile.scala 32:15]
  assign io_log_2 = regs__T_7_data; // @[RegFile.scala 32:15]
  assign io_log_3 = regs__T_8_data; // @[RegFile.scala 32:15]
  assign io_log_4 = regs__T_9_data; // @[RegFile.scala 32:15]
  assign io_log_5 = regs__T_10_data; // @[RegFile.scala 32:15]
  assign io_log_6 = regs__T_11_data; // @[RegFile.scala 32:15]
  assign io_log_7 = regs__T_12_data; // @[RegFile.scala 32:15]
  assign io_log_8 = regs__T_13_data; // @[RegFile.scala 32:15]
  assign io_log_9 = regs__T_14_data; // @[RegFile.scala 32:15]
  assign io_log_10 = regs__T_15_data; // @[RegFile.scala 32:15]
  assign io_log_11 = regs__T_16_data; // @[RegFile.scala 32:15]
  assign io_log_12 = regs__T_17_data; // @[RegFile.scala 32:15]
  assign io_log_13 = regs__T_18_data; // @[RegFile.scala 32:15]
  assign io_log_14 = regs__T_19_data; // @[RegFile.scala 32:15]
  assign io_log_15 = regs__T_20_data; // @[RegFile.scala 32:15]
  assign io_log_16 = regs__T_21_data; // @[RegFile.scala 32:15]
  assign io_log_17 = regs__T_22_data; // @[RegFile.scala 32:15]
  assign io_log_18 = regs__T_23_data; // @[RegFile.scala 32:15]
  assign io_log_19 = regs__T_24_data; // @[RegFile.scala 32:15]
  assign io_log_20 = regs__T_25_data; // @[RegFile.scala 32:15]
  assign io_log_21 = regs__T_26_data; // @[RegFile.scala 32:15]
  assign io_log_22 = regs__T_27_data; // @[RegFile.scala 32:15]
  assign io_log_23 = regs__T_28_data; // @[RegFile.scala 32:15]
  assign io_log_24 = regs__T_29_data; // @[RegFile.scala 32:15]
  assign io_log_25 = regs__T_30_data; // @[RegFile.scala 32:15]
  assign io_log_26 = regs__T_31_data; // @[RegFile.scala 32:15]
  assign io_log_27 = regs__T_32_data; // @[RegFile.scala 32:15]
  assign io_log_28 = regs__T_33_data; // @[RegFile.scala 32:15]
  assign io_log_29 = regs__T_34_data; // @[RegFile.scala 32:15]
  assign io_log_30 = regs__T_35_data; // @[RegFile.scala 32:15]
  assign io_log_31 = regs__T_36_data; // @[RegFile.scala 32:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(regs__T_en & regs__T_mask) begin
      regs[regs__T_addr] <= regs__T_data; // @[RegFile.scala 14:17]
    end
    if(regs__T_4_en & regs__T_4_mask) begin
      regs[regs__T_4_addr] <= regs__T_4_data; // @[RegFile.scala 14:17]
    end
  end
endmodule
module PTW(
  input         clock,
  input         reset,
  input  [9:0]  io_root_p2,
  input  [9:0]  io_root_p1,
  output        io_req_ready,
  input         io_req_valid,
  input  [9:0]  io_req_bits_p2,
  input  [9:0]  io_req_bits_p1,
  input         io_rsp_ready,
  output        io_rsp_valid,
  output [9:0]  io_rsp_bits_ppn_p2,
  output [9:0]  io_rsp_bits_ppn_p1,
  output        io_rsp_bits_U,
  output        io_rsp_bits_X,
  output        io_rsp_bits_W,
  output        io_rsp_bits_R,
  output        io_rsp_bits_V,
  output [31:0] io_mem_addr,
  output [3:0]  io_mem_mode,
  input  [31:0] io_mem_rdata,
  input         io_mem_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] status; // @[PTW.scala 53:23]
  reg [9:0] req_p1; // @[PTW.scala 54:23]
  wire  pte_V = io_mem_rdata[0]; // @[PTW.scala 55:37]
  wire  pte_R = io_mem_rdata[1]; // @[PTW.scala 55:37]
  wire  pte_W = io_mem_rdata[2]; // @[PTW.scala 55:37]
  wire  pte_X = io_mem_rdata[3]; // @[PTW.scala 55:37]
  wire  pte_U = io_mem_rdata[4]; // @[PTW.scala 55:37]
  wire [9:0] pte_ppn_p1 = io_mem_rdata[19:10]; // @[PTW.scala 55:37]
  wire [9:0] pte_ppn_p2 = io_mem_rdata[29:20]; // @[PTW.scala 55:37]
  wire  _T_16 = 2'h0 == status; // @[Conditional.scala 37:30]
  wire [11:0] _GEN_116 = {io_req_bits_p2, 2'h0}; // @[PTW.scala 72:54]
  wire [12:0] _T_17 = {{1'd0}, _GEN_116}; // @[PTW.scala 72:54]
  wire [31:0] _T_20 = {io_root_p2,io_root_p1,_T_17[11:0]}; // @[PTW.scala 12:53]
  wire [31:0] _GEN_1 = io_req_valid ? _T_20 : 32'h0; // @[PTW.scala 69:26]
  wire  _T_21 = 2'h1 == status; // @[Conditional.scala 37:30]
  wire  _T_22 = ~pte_V; // @[PTW.scala 80:14]
  wire  _T_23 = ~pte_R; // @[PTW.scala 35:26]
  wire  _T_24 = pte_V & _T_23; // @[PTW.scala 35:23]
  wire  _T_25 = ~pte_W; // @[PTW.scala 35:32]
  wire  _T_26 = _T_24 & _T_25; // @[PTW.scala 35:29]
  wire  _T_27 = ~_T_26; // @[PTW.scala 85:20]
  wire  _T_28 = |pte_ppn_p1; // @[PTW.scala 89:40]
  wire  _T_29 = ~_T_28; // @[PTW.scala 89:28]
  wire [11:0] _GEN_117 = {req_p1, 2'h0}; // @[PTW.scala 96:48]
  wire [12:0] _T_30 = {{1'd0}, _GEN_117}; // @[PTW.scala 96:48]
  wire [31:0] _T_33 = {pte_ppn_p2,pte_ppn_p1,_T_30[11:0]}; // @[PTW.scala 12:53]
  wire  _GEN_7 = _T_27 & _T_29; // @[PTW.scala 85:32]
  wire  _GEN_8 = _T_27 & pte_R; // @[PTW.scala 85:32]
  wire  _GEN_9 = _T_27 & pte_W; // @[PTW.scala 85:32]
  wire  _GEN_10 = _T_27 & pte_X; // @[PTW.scala 85:32]
  wire  _GEN_11 = _T_27 & pte_U; // @[PTW.scala 85:32]
  wire [9:0] _GEN_16 = _T_27 ? req_p1 : 10'h0; // @[PTW.scala 85:32]
  wire [9:0] _GEN_17 = _T_27 ? pte_ppn_p2 : 10'h0; // @[PTW.scala 85:32]
  wire  _GEN_20 = _T_27 ? 1'h0 : 1'h1; // @[PTW.scala 85:32]
  wire [31:0] _GEN_21 = _T_27 ? 32'h0 : _T_33; // @[PTW.scala 85:32]
  wire  _GEN_22 = _T_22 | _T_27; // @[PTW.scala 80:22]
  wire  _GEN_24 = _T_22 ? 1'h0 : _GEN_7; // @[PTW.scala 80:22]
  wire  _GEN_25 = _T_22 ? 1'h0 : _GEN_8; // @[PTW.scala 80:22]
  wire  _GEN_26 = _T_22 ? 1'h0 : _GEN_9; // @[PTW.scala 80:22]
  wire  _GEN_27 = _T_22 ? 1'h0 : _GEN_10; // @[PTW.scala 80:22]
  wire  _GEN_28 = _T_22 ? 1'h0 : _GEN_11; // @[PTW.scala 80:22]
  wire [9:0] _GEN_33 = _T_22 ? 10'h0 : _GEN_16; // @[PTW.scala 80:22]
  wire [9:0] _GEN_34 = _T_22 ? 10'h0 : _GEN_17; // @[PTW.scala 80:22]
  wire  _GEN_36 = _T_22 ? 1'h0 : _GEN_20; // @[PTW.scala 80:22]
  wire [31:0] _GEN_37 = _T_22 ? 32'h0 : _GEN_21; // @[PTW.scala 80:22]
  wire  _GEN_38 = io_mem_ok & _GEN_22; // @[PTW.scala 78:20]
  wire  _GEN_40 = io_mem_ok & _GEN_24; // @[PTW.scala 78:20]
  wire  _GEN_41 = io_mem_ok & _GEN_25; // @[PTW.scala 78:20]
  wire  _GEN_42 = io_mem_ok & _GEN_26; // @[PTW.scala 78:20]
  wire  _GEN_43 = io_mem_ok & _GEN_27; // @[PTW.scala 78:20]
  wire  _GEN_44 = io_mem_ok & _GEN_28; // @[PTW.scala 78:20]
  wire [9:0] _GEN_49 = io_mem_ok ? _GEN_33 : 10'h0; // @[PTW.scala 78:20]
  wire [9:0] _GEN_50 = io_mem_ok ? _GEN_34 : 10'h0; // @[PTW.scala 78:20]
  wire  _GEN_52 = io_mem_ok & _GEN_36; // @[PTW.scala 78:20]
  wire [31:0] _GEN_53 = io_mem_ok ? _GEN_37 : 32'h0; // @[PTW.scala 78:20]
  wire  _T_34 = 2'h2 == status; // @[Conditional.scala 37:30]
  wire  _T_35 = pte_R | pte_W; // @[PTW.scala 36:30]
  wire  _T_36 = pte_V & _T_35; // @[PTW.scala 36:24]
  wire  _GEN_55 = io_mem_ok & _T_36; // @[PTW.scala 102:20]
  wire  _GEN_56 = io_mem_ok & pte_R; // @[PTW.scala 102:20]
  wire  _GEN_57 = io_mem_ok & pte_W; // @[PTW.scala 102:20]
  wire  _GEN_58 = io_mem_ok & pte_X; // @[PTW.scala 102:20]
  wire  _GEN_59 = io_mem_ok & pte_U; // @[PTW.scala 102:20]
  wire [9:0] _GEN_64 = io_mem_ok ? pte_ppn_p1 : 10'h0; // @[PTW.scala 102:20]
  wire [9:0] _GEN_65 = io_mem_ok ? pte_ppn_p2 : 10'h0; // @[PTW.scala 102:20]
  wire  _GEN_68 = _T_34 & io_mem_ok; // @[Conditional.scala 39:67]
  wire  _GEN_69 = _T_34 & _GEN_55; // @[Conditional.scala 39:67]
  wire  _GEN_70 = _T_34 & _GEN_56; // @[Conditional.scala 39:67]
  wire  _GEN_71 = _T_34 & _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_72 = _T_34 & _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_73 = _T_34 & _GEN_59; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_78 = _T_34 ? _GEN_64 : 10'h0; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_79 = _T_34 ? _GEN_65 : 10'h0; // @[Conditional.scala 39:67]
  wire  _GEN_82 = _T_21 ? _GEN_38 : _GEN_68; // @[Conditional.scala 39:67]
  wire  _GEN_84 = _T_21 ? _GEN_40 : _GEN_69; // @[Conditional.scala 39:67]
  wire  _GEN_85 = _T_21 ? _GEN_41 : _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_86 = _T_21 ? _GEN_42 : _GEN_71; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_21 ? _GEN_43 : _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_88 = _T_21 ? _GEN_44 : _GEN_73; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_93 = _T_21 ? _GEN_49 : _GEN_78; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_94 = _T_21 ? _GEN_50 : _GEN_79; // @[Conditional.scala 39:67]
  wire  _GEN_96 = _T_21 & _GEN_52; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_97 = _T_21 ? _GEN_53 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_98 = _T_16 ? io_req_valid : _GEN_96; // @[Conditional.scala 40:58]
  assign io_req_ready = status == 2'h0; // @[PTW.scala 58:16]
  assign io_rsp_valid = _T_16 ? 1'h0 : _GEN_82; // @[PTW.scala 64:16 PTW.scala 81:24 PTW.scala 86:24 PTW.scala 103:22]
  assign io_rsp_bits_ppn_p2 = _T_16 ? 10'h0 : _GEN_94; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 104:21]
  assign io_rsp_bits_ppn_p1 = _T_16 ? 10'h0 : _GEN_93; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 88:30 PTW.scala 104:21]
  assign io_rsp_bits_U = _T_16 ? 1'h0 : _GEN_88; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 104:21]
  assign io_rsp_bits_X = _T_16 ? 1'h0 : _GEN_87; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 104:21]
  assign io_rsp_bits_W = _T_16 ? 1'h0 : _GEN_86; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 104:21]
  assign io_rsp_bits_R = _T_16 ? 1'h0 : _GEN_85; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 104:21]
  assign io_rsp_bits_V = _T_16 ? 1'h0 : _GEN_84; // @[PTW.scala 65:15 PTW.scala 87:23 PTW.scala 89:25 PTW.scala 104:21 PTW.scala 105:23]
  assign io_mem_addr = _T_16 ? _GEN_1 : _GEN_97; // @[PTW.scala 62:15 PTW.scala 72:21 PTW.scala 96:23]
  assign io_mem_mode = {{3'd0}, _GEN_98}; // @[PTW.scala 61:15 PTW.scala 71:21 PTW.scala 95:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  status = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  req_p1 = _RAND_1[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      status <= 2'h0;
    end else if (_T_16) begin
      if (io_req_valid) begin
        status <= 2'h1;
      end
    end else if (_T_21) begin
      if (io_mem_ok) begin
        if (_T_22) begin
          if (io_rsp_ready) begin
            status <= 2'h0;
          end
        end else if (_T_27) begin
          if (io_rsp_ready) begin
            status <= 2'h0;
          end
        end else begin
          status <= 2'h2;
        end
      end
    end else if (_T_34) begin
      if (io_mem_ok) begin
        if (io_rsp_ready) begin
          status <= 2'h0;
        end
      end
    end
    if (reset) begin
      req_p1 <= 10'h0;
    end else if (_T_16) begin
      if (io_req_valid) begin
        req_p1 <= io_req_bits_p1;
      end
    end
  end
endmodule
module TLB(
  input        clock,
  input        reset,
  input        io_query_req_valid,
  input  [9:0] io_query_req_bits_p2,
  input  [9:0] io_query_req_bits_p1,
  output       io_query_rsp_valid,
  output [9:0] io_query_rsp_bits_ppn_p2,
  output [9:0] io_query_rsp_bits_ppn_p1,
  output       io_query_rsp_bits_U,
  output       io_query_rsp_bits_X,
  output       io_query_rsp_bits_V,
  input        io_query2_req_valid,
  input  [9:0] io_query2_req_bits_p2,
  input  [9:0] io_query2_req_bits_p1,
  output       io_query2_rsp_valid,
  output [9:0] io_query2_rsp_bits_ppn_p2,
  output [9:0] io_query2_rsp_bits_ppn_p1,
  output       io_query2_rsp_bits_U,
  output       io_query2_rsp_bits_X,
  output       io_query2_rsp_bits_W,
  output       io_query2_rsp_bits_R,
  output       io_query2_rsp_bits_V,
  input  [1:0] io_modify_mode,
  input  [9:0] io_modify_vpn_p2,
  input  [9:0] io_modify_vpn_p1,
  input  [9:0] io_modify_pte_ppn_p2,
  input  [9:0] io_modify_pte_ppn_p1,
  input        io_modify_pte_U,
  input        io_modify_pte_X,
  input        io_modify_pte_W,
  input        io_modify_pte_R,
  input        io_modify_pte_V
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
  reg  entries_valid [0:31]; // @[TLB.scala 38:20]
  wire  entries_valid__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_3_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_4_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_5_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_6_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_7_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_8_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_9_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_10_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_11_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_12_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_13_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_14_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_15_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_16_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_17_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_18_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_19_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_20_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_21_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_22_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_23_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_24_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_25_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_26_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_27_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_28_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_29_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_30_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_31_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_32_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_33_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_34_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_57_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_58_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_59_en; // @[TLB.scala 38:20]
  wire  entries_valid__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_valid__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_valid__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_valid__T_65_en; // @[TLB.scala 38:20]
  reg [9:0] entries_vpn_p2 [0:31]; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_39_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_49_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_61_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_3_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_4_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_5_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_6_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_7_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_8_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_9_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_10_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_11_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_12_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_13_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_14_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_15_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_16_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_17_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_18_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_19_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_20_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_21_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_22_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_23_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_24_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_25_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_26_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_27_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_28_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_29_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_30_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_31_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_32_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_33_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_34_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_57_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_58_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_59_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p2__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p2__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p2__T_65_en; // @[TLB.scala 38:20]
  reg [9:0] entries_vpn_p1 [0:31]; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_39_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_49_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_61_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_3_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_4_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_5_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_6_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_7_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_8_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_9_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_10_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_11_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_12_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_13_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_14_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_15_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_16_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_17_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_18_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_19_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_20_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_21_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_22_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_23_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_24_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_25_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_26_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_27_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_28_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_29_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_30_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_31_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_32_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_33_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_34_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_57_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_58_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_59_en; // @[TLB.scala 38:20]
  wire [9:0] entries_vpn_p1__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_vpn_p1__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_vpn_p1__T_65_en; // @[TLB.scala 38:20]
  reg [9:0] entries_pte_ppn_p2 [0:31]; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_39_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_49_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_61_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_3_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_4_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_5_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_6_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_7_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_8_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_9_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_10_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_11_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_12_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_13_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_14_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_15_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_16_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_17_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_18_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_19_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_20_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_21_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_22_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_23_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_24_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_25_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_26_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_27_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_28_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_29_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_30_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_31_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_32_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_33_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_34_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_57_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_58_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_59_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p2__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p2__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p2__T_65_en; // @[TLB.scala 38:20]
  reg [9:0] entries_pte_ppn_p1 [0:31]; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_39_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_49_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_61_addr; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_3_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_4_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_5_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_6_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_7_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_8_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_9_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_10_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_11_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_12_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_13_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_14_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_15_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_16_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_17_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_18_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_19_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_20_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_21_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_22_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_23_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_24_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_25_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_26_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_27_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_28_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_29_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_30_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_31_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_32_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_33_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_34_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_57_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_58_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_59_en; // @[TLB.scala 38:20]
  wire [9:0] entries_pte_ppn_p1__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_ppn_p1__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_ppn_p1__T_65_en; // @[TLB.scala 38:20]
  reg  entries_pte_U [0:31]; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_3_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_4_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_5_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_6_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_7_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_8_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_9_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_10_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_11_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_12_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_13_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_14_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_15_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_16_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_17_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_18_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_19_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_20_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_21_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_22_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_23_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_24_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_25_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_26_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_27_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_28_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_29_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_30_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_31_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_32_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_33_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_34_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_57_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_58_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_59_en; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_U__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_U__T_65_en; // @[TLB.scala 38:20]
  reg  entries_pte_X [0:31]; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_3_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_4_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_5_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_6_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_7_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_8_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_9_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_10_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_11_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_12_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_13_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_14_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_15_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_16_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_17_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_18_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_19_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_20_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_21_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_22_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_23_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_24_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_25_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_26_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_27_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_28_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_29_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_30_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_31_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_32_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_33_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_34_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_57_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_58_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_59_en; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_X__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_X__T_65_en; // @[TLB.scala 38:20]
  reg  entries_pte_W [0:31]; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_3_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_4_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_5_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_6_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_7_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_8_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_9_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_10_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_11_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_12_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_13_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_14_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_15_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_16_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_17_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_18_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_19_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_20_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_21_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_22_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_23_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_24_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_25_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_26_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_27_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_28_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_29_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_30_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_31_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_32_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_33_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_34_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_57_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_58_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_59_en; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_W__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_W__T_65_en; // @[TLB.scala 38:20]
  reg  entries_pte_R [0:31]; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_3_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_4_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_5_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_6_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_7_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_8_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_9_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_10_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_11_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_12_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_13_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_14_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_15_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_16_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_17_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_18_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_19_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_20_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_21_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_22_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_23_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_24_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_25_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_26_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_27_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_28_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_29_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_30_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_31_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_32_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_33_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_34_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_57_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_58_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_59_en; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_R__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_R__T_65_en; // @[TLB.scala 38:20]
  reg  entries_pte_V [0:31]; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_39_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_39_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_49_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_49_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_61_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_61_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_3_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_3_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_3_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_3_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_4_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_4_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_4_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_4_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_5_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_5_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_5_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_5_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_6_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_6_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_6_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_6_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_7_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_7_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_7_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_7_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_8_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_8_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_8_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_8_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_9_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_9_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_9_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_9_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_10_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_10_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_10_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_10_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_11_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_11_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_11_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_11_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_12_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_12_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_12_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_12_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_13_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_13_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_13_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_13_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_14_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_14_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_14_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_14_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_15_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_15_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_15_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_15_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_16_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_16_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_16_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_16_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_17_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_17_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_17_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_17_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_18_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_18_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_18_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_18_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_19_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_19_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_19_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_19_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_20_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_20_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_20_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_20_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_21_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_21_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_21_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_21_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_22_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_22_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_22_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_22_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_23_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_23_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_23_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_23_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_24_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_24_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_24_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_24_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_25_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_25_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_25_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_25_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_26_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_26_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_26_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_26_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_27_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_27_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_27_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_27_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_28_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_28_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_28_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_28_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_29_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_29_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_29_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_29_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_30_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_30_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_30_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_30_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_31_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_31_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_31_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_31_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_32_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_32_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_32_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_32_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_33_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_33_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_33_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_33_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_34_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_34_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_34_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_34_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_57_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_57_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_57_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_57_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_58_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_58_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_58_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_58_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_59_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_59_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_59_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_59_en; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_65_data; // @[TLB.scala 38:20]
  wire [4:0] entries_pte_V__T_65_addr; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_65_mask; // @[TLB.scala 38:20]
  wire  entries_pte_V__T_65_en; // @[TLB.scala 38:20]
  wire  _T_1 = io_modify_mode == 2'h3; // @[TLB.scala 45:39]
  wire [9:0] _T_37 = io_query_req_bits_p2 ^ io_query_req_bits_p1; // @[TLB.scala 51:34]
  wire  _T_40 = io_query_req_valid & entries_valid__T_39_data; // @[TLB.scala 67:34]
  wire [19:0] _T_41 = {entries_vpn_p2__T_39_data,entries_vpn_p1__T_39_data}; // @[TLB.scala 67:62]
  wire [19:0] _T_42 = {io_query_req_bits_p2,io_query_req_bits_p1}; // @[TLB.scala 67:84]
  wire  _T_43 = _T_41 == _T_42; // @[TLB.scala 67:69]
  wire  _T_44 = _T_40 & _T_43; // @[TLB.scala 67:49]
  wire [9:0] _T_47 = io_query2_req_bits_p2 ^ io_query2_req_bits_p1; // @[TLB.scala 51:34]
  wire  _T_50 = io_query2_req_valid & entries_valid__T_49_data; // @[TLB.scala 67:34]
  wire [19:0] _T_51 = {entries_vpn_p2__T_49_data,entries_vpn_p1__T_49_data}; // @[TLB.scala 67:62]
  wire [19:0] _T_52 = {io_query2_req_bits_p2,io_query2_req_bits_p1}; // @[TLB.scala 67:84]
  wire  _T_53 = _T_51 == _T_52; // @[TLB.scala 67:69]
  wire  _T_54 = _T_50 & _T_53; // @[TLB.scala 67:49]
  wire [9:0] _T_55 = io_modify_vpn_p2 ^ io_modify_vpn_p1; // @[TLB.scala 51:34]
  wire  _T_60 = io_modify_mode == 2'h2; // @[TLB.scala 88:23]
  wire [19:0] _T_62 = {entries_vpn_p2__T_61_data,entries_vpn_p1__T_61_data}; // @[TLB.scala 89:26]
  wire [19:0] _T_63 = {io_modify_vpn_p2,io_modify_vpn_p1}; // @[TLB.scala 89:51]
  wire  _T_64 = _T_62 == _T_63; // @[TLB.scala 89:33]
  assign entries_valid__T_39_addr = _T_37[4:0];
  assign entries_valid__T_39_data = entries_valid[entries_valid__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_valid__T_49_addr = _T_47[4:0];
  assign entries_valid__T_49_data = entries_valid[entries_valid__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_valid__T_61_addr = _T_55[4:0];
  assign entries_valid__T_61_data = entries_valid[entries_valid__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_valid__T_3_data = 1'h0;
  assign entries_valid__T_3_addr = 5'h0;
  assign entries_valid__T_3_mask = 1'h1;
  assign entries_valid__T_3_en = reset | _T_1;
  assign entries_valid__T_4_data = 1'h0;
  assign entries_valid__T_4_addr = 5'h1;
  assign entries_valid__T_4_mask = 1'h1;
  assign entries_valid__T_4_en = reset | _T_1;
  assign entries_valid__T_5_data = 1'h0;
  assign entries_valid__T_5_addr = 5'h2;
  assign entries_valid__T_5_mask = 1'h1;
  assign entries_valid__T_5_en = reset | _T_1;
  assign entries_valid__T_6_data = 1'h0;
  assign entries_valid__T_6_addr = 5'h3;
  assign entries_valid__T_6_mask = 1'h1;
  assign entries_valid__T_6_en = reset | _T_1;
  assign entries_valid__T_7_data = 1'h0;
  assign entries_valid__T_7_addr = 5'h4;
  assign entries_valid__T_7_mask = 1'h1;
  assign entries_valid__T_7_en = reset | _T_1;
  assign entries_valid__T_8_data = 1'h0;
  assign entries_valid__T_8_addr = 5'h5;
  assign entries_valid__T_8_mask = 1'h1;
  assign entries_valid__T_8_en = reset | _T_1;
  assign entries_valid__T_9_data = 1'h0;
  assign entries_valid__T_9_addr = 5'h6;
  assign entries_valid__T_9_mask = 1'h1;
  assign entries_valid__T_9_en = reset | _T_1;
  assign entries_valid__T_10_data = 1'h0;
  assign entries_valid__T_10_addr = 5'h7;
  assign entries_valid__T_10_mask = 1'h1;
  assign entries_valid__T_10_en = reset | _T_1;
  assign entries_valid__T_11_data = 1'h0;
  assign entries_valid__T_11_addr = 5'h8;
  assign entries_valid__T_11_mask = 1'h1;
  assign entries_valid__T_11_en = reset | _T_1;
  assign entries_valid__T_12_data = 1'h0;
  assign entries_valid__T_12_addr = 5'h9;
  assign entries_valid__T_12_mask = 1'h1;
  assign entries_valid__T_12_en = reset | _T_1;
  assign entries_valid__T_13_data = 1'h0;
  assign entries_valid__T_13_addr = 5'ha;
  assign entries_valid__T_13_mask = 1'h1;
  assign entries_valid__T_13_en = reset | _T_1;
  assign entries_valid__T_14_data = 1'h0;
  assign entries_valid__T_14_addr = 5'hb;
  assign entries_valid__T_14_mask = 1'h1;
  assign entries_valid__T_14_en = reset | _T_1;
  assign entries_valid__T_15_data = 1'h0;
  assign entries_valid__T_15_addr = 5'hc;
  assign entries_valid__T_15_mask = 1'h1;
  assign entries_valid__T_15_en = reset | _T_1;
  assign entries_valid__T_16_data = 1'h0;
  assign entries_valid__T_16_addr = 5'hd;
  assign entries_valid__T_16_mask = 1'h1;
  assign entries_valid__T_16_en = reset | _T_1;
  assign entries_valid__T_17_data = 1'h0;
  assign entries_valid__T_17_addr = 5'he;
  assign entries_valid__T_17_mask = 1'h1;
  assign entries_valid__T_17_en = reset | _T_1;
  assign entries_valid__T_18_data = 1'h0;
  assign entries_valid__T_18_addr = 5'hf;
  assign entries_valid__T_18_mask = 1'h1;
  assign entries_valid__T_18_en = reset | _T_1;
  assign entries_valid__T_19_data = 1'h0;
  assign entries_valid__T_19_addr = 5'h10;
  assign entries_valid__T_19_mask = 1'h1;
  assign entries_valid__T_19_en = reset | _T_1;
  assign entries_valid__T_20_data = 1'h0;
  assign entries_valid__T_20_addr = 5'h11;
  assign entries_valid__T_20_mask = 1'h1;
  assign entries_valid__T_20_en = reset | _T_1;
  assign entries_valid__T_21_data = 1'h0;
  assign entries_valid__T_21_addr = 5'h12;
  assign entries_valid__T_21_mask = 1'h1;
  assign entries_valid__T_21_en = reset | _T_1;
  assign entries_valid__T_22_data = 1'h0;
  assign entries_valid__T_22_addr = 5'h13;
  assign entries_valid__T_22_mask = 1'h1;
  assign entries_valid__T_22_en = reset | _T_1;
  assign entries_valid__T_23_data = 1'h0;
  assign entries_valid__T_23_addr = 5'h14;
  assign entries_valid__T_23_mask = 1'h1;
  assign entries_valid__T_23_en = reset | _T_1;
  assign entries_valid__T_24_data = 1'h0;
  assign entries_valid__T_24_addr = 5'h15;
  assign entries_valid__T_24_mask = 1'h1;
  assign entries_valid__T_24_en = reset | _T_1;
  assign entries_valid__T_25_data = 1'h0;
  assign entries_valid__T_25_addr = 5'h16;
  assign entries_valid__T_25_mask = 1'h1;
  assign entries_valid__T_25_en = reset | _T_1;
  assign entries_valid__T_26_data = 1'h0;
  assign entries_valid__T_26_addr = 5'h17;
  assign entries_valid__T_26_mask = 1'h1;
  assign entries_valid__T_26_en = reset | _T_1;
  assign entries_valid__T_27_data = 1'h0;
  assign entries_valid__T_27_addr = 5'h18;
  assign entries_valid__T_27_mask = 1'h1;
  assign entries_valid__T_27_en = reset | _T_1;
  assign entries_valid__T_28_data = 1'h0;
  assign entries_valid__T_28_addr = 5'h19;
  assign entries_valid__T_28_mask = 1'h1;
  assign entries_valid__T_28_en = reset | _T_1;
  assign entries_valid__T_29_data = 1'h0;
  assign entries_valid__T_29_addr = 5'h1a;
  assign entries_valid__T_29_mask = 1'h1;
  assign entries_valid__T_29_en = reset | _T_1;
  assign entries_valid__T_30_data = 1'h0;
  assign entries_valid__T_30_addr = 5'h1b;
  assign entries_valid__T_30_mask = 1'h1;
  assign entries_valid__T_30_en = reset | _T_1;
  assign entries_valid__T_31_data = 1'h0;
  assign entries_valid__T_31_addr = 5'h1c;
  assign entries_valid__T_31_mask = 1'h1;
  assign entries_valid__T_31_en = reset | _T_1;
  assign entries_valid__T_32_data = 1'h0;
  assign entries_valid__T_32_addr = 5'h1d;
  assign entries_valid__T_32_mask = 1'h1;
  assign entries_valid__T_32_en = reset | _T_1;
  assign entries_valid__T_33_data = 1'h0;
  assign entries_valid__T_33_addr = 5'h1e;
  assign entries_valid__T_33_mask = 1'h1;
  assign entries_valid__T_33_en = reset | _T_1;
  assign entries_valid__T_34_data = 1'h0;
  assign entries_valid__T_34_addr = 5'h1f;
  assign entries_valid__T_34_mask = 1'h1;
  assign entries_valid__T_34_en = reset | _T_1;
  assign entries_valid__T_57_data = 1'h1;
  assign entries_valid__T_57_addr = _T_55[4:0];
  assign entries_valid__T_57_mask = 1'h1;
  assign entries_valid__T_57_en = io_modify_mode == 2'h1;
  assign entries_valid__T_58_data = 1'h0;
  assign entries_valid__T_58_addr = _T_55[4:0];
  assign entries_valid__T_58_mask = 1'h0;
  assign entries_valid__T_58_en = io_modify_mode == 2'h1;
  assign entries_valid__T_59_data = 1'h0;
  assign entries_valid__T_59_addr = _T_55[4:0];
  assign entries_valid__T_59_mask = 1'h0;
  assign entries_valid__T_59_en = io_modify_mode == 2'h1;
  assign entries_valid__T_65_data = 1'h0;
  assign entries_valid__T_65_addr = _T_55[4:0];
  assign entries_valid__T_65_mask = 1'h1;
  assign entries_valid__T_65_en = _T_60 & _T_64;
  assign entries_vpn_p2__T_39_addr = _T_37[4:0];
  assign entries_vpn_p2__T_39_data = entries_vpn_p2[entries_vpn_p2__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p2__T_49_addr = _T_47[4:0];
  assign entries_vpn_p2__T_49_data = entries_vpn_p2[entries_vpn_p2__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p2__T_61_addr = _T_55[4:0];
  assign entries_vpn_p2__T_61_data = entries_vpn_p2[entries_vpn_p2__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p2__T_3_data = 10'h0;
  assign entries_vpn_p2__T_3_addr = 5'h0;
  assign entries_vpn_p2__T_3_mask = 1'h0;
  assign entries_vpn_p2__T_3_en = reset | _T_1;
  assign entries_vpn_p2__T_4_data = 10'h0;
  assign entries_vpn_p2__T_4_addr = 5'h1;
  assign entries_vpn_p2__T_4_mask = 1'h0;
  assign entries_vpn_p2__T_4_en = reset | _T_1;
  assign entries_vpn_p2__T_5_data = 10'h0;
  assign entries_vpn_p2__T_5_addr = 5'h2;
  assign entries_vpn_p2__T_5_mask = 1'h0;
  assign entries_vpn_p2__T_5_en = reset | _T_1;
  assign entries_vpn_p2__T_6_data = 10'h0;
  assign entries_vpn_p2__T_6_addr = 5'h3;
  assign entries_vpn_p2__T_6_mask = 1'h0;
  assign entries_vpn_p2__T_6_en = reset | _T_1;
  assign entries_vpn_p2__T_7_data = 10'h0;
  assign entries_vpn_p2__T_7_addr = 5'h4;
  assign entries_vpn_p2__T_7_mask = 1'h0;
  assign entries_vpn_p2__T_7_en = reset | _T_1;
  assign entries_vpn_p2__T_8_data = 10'h0;
  assign entries_vpn_p2__T_8_addr = 5'h5;
  assign entries_vpn_p2__T_8_mask = 1'h0;
  assign entries_vpn_p2__T_8_en = reset | _T_1;
  assign entries_vpn_p2__T_9_data = 10'h0;
  assign entries_vpn_p2__T_9_addr = 5'h6;
  assign entries_vpn_p2__T_9_mask = 1'h0;
  assign entries_vpn_p2__T_9_en = reset | _T_1;
  assign entries_vpn_p2__T_10_data = 10'h0;
  assign entries_vpn_p2__T_10_addr = 5'h7;
  assign entries_vpn_p2__T_10_mask = 1'h0;
  assign entries_vpn_p2__T_10_en = reset | _T_1;
  assign entries_vpn_p2__T_11_data = 10'h0;
  assign entries_vpn_p2__T_11_addr = 5'h8;
  assign entries_vpn_p2__T_11_mask = 1'h0;
  assign entries_vpn_p2__T_11_en = reset | _T_1;
  assign entries_vpn_p2__T_12_data = 10'h0;
  assign entries_vpn_p2__T_12_addr = 5'h9;
  assign entries_vpn_p2__T_12_mask = 1'h0;
  assign entries_vpn_p2__T_12_en = reset | _T_1;
  assign entries_vpn_p2__T_13_data = 10'h0;
  assign entries_vpn_p2__T_13_addr = 5'ha;
  assign entries_vpn_p2__T_13_mask = 1'h0;
  assign entries_vpn_p2__T_13_en = reset | _T_1;
  assign entries_vpn_p2__T_14_data = 10'h0;
  assign entries_vpn_p2__T_14_addr = 5'hb;
  assign entries_vpn_p2__T_14_mask = 1'h0;
  assign entries_vpn_p2__T_14_en = reset | _T_1;
  assign entries_vpn_p2__T_15_data = 10'h0;
  assign entries_vpn_p2__T_15_addr = 5'hc;
  assign entries_vpn_p2__T_15_mask = 1'h0;
  assign entries_vpn_p2__T_15_en = reset | _T_1;
  assign entries_vpn_p2__T_16_data = 10'h0;
  assign entries_vpn_p2__T_16_addr = 5'hd;
  assign entries_vpn_p2__T_16_mask = 1'h0;
  assign entries_vpn_p2__T_16_en = reset | _T_1;
  assign entries_vpn_p2__T_17_data = 10'h0;
  assign entries_vpn_p2__T_17_addr = 5'he;
  assign entries_vpn_p2__T_17_mask = 1'h0;
  assign entries_vpn_p2__T_17_en = reset | _T_1;
  assign entries_vpn_p2__T_18_data = 10'h0;
  assign entries_vpn_p2__T_18_addr = 5'hf;
  assign entries_vpn_p2__T_18_mask = 1'h0;
  assign entries_vpn_p2__T_18_en = reset | _T_1;
  assign entries_vpn_p2__T_19_data = 10'h0;
  assign entries_vpn_p2__T_19_addr = 5'h10;
  assign entries_vpn_p2__T_19_mask = 1'h0;
  assign entries_vpn_p2__T_19_en = reset | _T_1;
  assign entries_vpn_p2__T_20_data = 10'h0;
  assign entries_vpn_p2__T_20_addr = 5'h11;
  assign entries_vpn_p2__T_20_mask = 1'h0;
  assign entries_vpn_p2__T_20_en = reset | _T_1;
  assign entries_vpn_p2__T_21_data = 10'h0;
  assign entries_vpn_p2__T_21_addr = 5'h12;
  assign entries_vpn_p2__T_21_mask = 1'h0;
  assign entries_vpn_p2__T_21_en = reset | _T_1;
  assign entries_vpn_p2__T_22_data = 10'h0;
  assign entries_vpn_p2__T_22_addr = 5'h13;
  assign entries_vpn_p2__T_22_mask = 1'h0;
  assign entries_vpn_p2__T_22_en = reset | _T_1;
  assign entries_vpn_p2__T_23_data = 10'h0;
  assign entries_vpn_p2__T_23_addr = 5'h14;
  assign entries_vpn_p2__T_23_mask = 1'h0;
  assign entries_vpn_p2__T_23_en = reset | _T_1;
  assign entries_vpn_p2__T_24_data = 10'h0;
  assign entries_vpn_p2__T_24_addr = 5'h15;
  assign entries_vpn_p2__T_24_mask = 1'h0;
  assign entries_vpn_p2__T_24_en = reset | _T_1;
  assign entries_vpn_p2__T_25_data = 10'h0;
  assign entries_vpn_p2__T_25_addr = 5'h16;
  assign entries_vpn_p2__T_25_mask = 1'h0;
  assign entries_vpn_p2__T_25_en = reset | _T_1;
  assign entries_vpn_p2__T_26_data = 10'h0;
  assign entries_vpn_p2__T_26_addr = 5'h17;
  assign entries_vpn_p2__T_26_mask = 1'h0;
  assign entries_vpn_p2__T_26_en = reset | _T_1;
  assign entries_vpn_p2__T_27_data = 10'h0;
  assign entries_vpn_p2__T_27_addr = 5'h18;
  assign entries_vpn_p2__T_27_mask = 1'h0;
  assign entries_vpn_p2__T_27_en = reset | _T_1;
  assign entries_vpn_p2__T_28_data = 10'h0;
  assign entries_vpn_p2__T_28_addr = 5'h19;
  assign entries_vpn_p2__T_28_mask = 1'h0;
  assign entries_vpn_p2__T_28_en = reset | _T_1;
  assign entries_vpn_p2__T_29_data = 10'h0;
  assign entries_vpn_p2__T_29_addr = 5'h1a;
  assign entries_vpn_p2__T_29_mask = 1'h0;
  assign entries_vpn_p2__T_29_en = reset | _T_1;
  assign entries_vpn_p2__T_30_data = 10'h0;
  assign entries_vpn_p2__T_30_addr = 5'h1b;
  assign entries_vpn_p2__T_30_mask = 1'h0;
  assign entries_vpn_p2__T_30_en = reset | _T_1;
  assign entries_vpn_p2__T_31_data = 10'h0;
  assign entries_vpn_p2__T_31_addr = 5'h1c;
  assign entries_vpn_p2__T_31_mask = 1'h0;
  assign entries_vpn_p2__T_31_en = reset | _T_1;
  assign entries_vpn_p2__T_32_data = 10'h0;
  assign entries_vpn_p2__T_32_addr = 5'h1d;
  assign entries_vpn_p2__T_32_mask = 1'h0;
  assign entries_vpn_p2__T_32_en = reset | _T_1;
  assign entries_vpn_p2__T_33_data = 10'h0;
  assign entries_vpn_p2__T_33_addr = 5'h1e;
  assign entries_vpn_p2__T_33_mask = 1'h0;
  assign entries_vpn_p2__T_33_en = reset | _T_1;
  assign entries_vpn_p2__T_34_data = 10'h0;
  assign entries_vpn_p2__T_34_addr = 5'h1f;
  assign entries_vpn_p2__T_34_mask = 1'h0;
  assign entries_vpn_p2__T_34_en = reset | _T_1;
  assign entries_vpn_p2__T_57_data = 10'h0;
  assign entries_vpn_p2__T_57_addr = _T_55[4:0];
  assign entries_vpn_p2__T_57_mask = 1'h0;
  assign entries_vpn_p2__T_57_en = io_modify_mode == 2'h1;
  assign entries_vpn_p2__T_58_data = io_modify_vpn_p2;
  assign entries_vpn_p2__T_58_addr = _T_55[4:0];
  assign entries_vpn_p2__T_58_mask = 1'h1;
  assign entries_vpn_p2__T_58_en = io_modify_mode == 2'h1;
  assign entries_vpn_p2__T_59_data = 10'h0;
  assign entries_vpn_p2__T_59_addr = _T_55[4:0];
  assign entries_vpn_p2__T_59_mask = 1'h0;
  assign entries_vpn_p2__T_59_en = io_modify_mode == 2'h1;
  assign entries_vpn_p2__T_65_data = 10'h0;
  assign entries_vpn_p2__T_65_addr = _T_55[4:0];
  assign entries_vpn_p2__T_65_mask = 1'h0;
  assign entries_vpn_p2__T_65_en = _T_60 & _T_64;
  assign entries_vpn_p1__T_39_addr = _T_37[4:0];
  assign entries_vpn_p1__T_39_data = entries_vpn_p1[entries_vpn_p1__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p1__T_49_addr = _T_47[4:0];
  assign entries_vpn_p1__T_49_data = entries_vpn_p1[entries_vpn_p1__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p1__T_61_addr = _T_55[4:0];
  assign entries_vpn_p1__T_61_data = entries_vpn_p1[entries_vpn_p1__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_vpn_p1__T_3_data = 10'h0;
  assign entries_vpn_p1__T_3_addr = 5'h0;
  assign entries_vpn_p1__T_3_mask = 1'h0;
  assign entries_vpn_p1__T_3_en = reset | _T_1;
  assign entries_vpn_p1__T_4_data = 10'h0;
  assign entries_vpn_p1__T_4_addr = 5'h1;
  assign entries_vpn_p1__T_4_mask = 1'h0;
  assign entries_vpn_p1__T_4_en = reset | _T_1;
  assign entries_vpn_p1__T_5_data = 10'h0;
  assign entries_vpn_p1__T_5_addr = 5'h2;
  assign entries_vpn_p1__T_5_mask = 1'h0;
  assign entries_vpn_p1__T_5_en = reset | _T_1;
  assign entries_vpn_p1__T_6_data = 10'h0;
  assign entries_vpn_p1__T_6_addr = 5'h3;
  assign entries_vpn_p1__T_6_mask = 1'h0;
  assign entries_vpn_p1__T_6_en = reset | _T_1;
  assign entries_vpn_p1__T_7_data = 10'h0;
  assign entries_vpn_p1__T_7_addr = 5'h4;
  assign entries_vpn_p1__T_7_mask = 1'h0;
  assign entries_vpn_p1__T_7_en = reset | _T_1;
  assign entries_vpn_p1__T_8_data = 10'h0;
  assign entries_vpn_p1__T_8_addr = 5'h5;
  assign entries_vpn_p1__T_8_mask = 1'h0;
  assign entries_vpn_p1__T_8_en = reset | _T_1;
  assign entries_vpn_p1__T_9_data = 10'h0;
  assign entries_vpn_p1__T_9_addr = 5'h6;
  assign entries_vpn_p1__T_9_mask = 1'h0;
  assign entries_vpn_p1__T_9_en = reset | _T_1;
  assign entries_vpn_p1__T_10_data = 10'h0;
  assign entries_vpn_p1__T_10_addr = 5'h7;
  assign entries_vpn_p1__T_10_mask = 1'h0;
  assign entries_vpn_p1__T_10_en = reset | _T_1;
  assign entries_vpn_p1__T_11_data = 10'h0;
  assign entries_vpn_p1__T_11_addr = 5'h8;
  assign entries_vpn_p1__T_11_mask = 1'h0;
  assign entries_vpn_p1__T_11_en = reset | _T_1;
  assign entries_vpn_p1__T_12_data = 10'h0;
  assign entries_vpn_p1__T_12_addr = 5'h9;
  assign entries_vpn_p1__T_12_mask = 1'h0;
  assign entries_vpn_p1__T_12_en = reset | _T_1;
  assign entries_vpn_p1__T_13_data = 10'h0;
  assign entries_vpn_p1__T_13_addr = 5'ha;
  assign entries_vpn_p1__T_13_mask = 1'h0;
  assign entries_vpn_p1__T_13_en = reset | _T_1;
  assign entries_vpn_p1__T_14_data = 10'h0;
  assign entries_vpn_p1__T_14_addr = 5'hb;
  assign entries_vpn_p1__T_14_mask = 1'h0;
  assign entries_vpn_p1__T_14_en = reset | _T_1;
  assign entries_vpn_p1__T_15_data = 10'h0;
  assign entries_vpn_p1__T_15_addr = 5'hc;
  assign entries_vpn_p1__T_15_mask = 1'h0;
  assign entries_vpn_p1__T_15_en = reset | _T_1;
  assign entries_vpn_p1__T_16_data = 10'h0;
  assign entries_vpn_p1__T_16_addr = 5'hd;
  assign entries_vpn_p1__T_16_mask = 1'h0;
  assign entries_vpn_p1__T_16_en = reset | _T_1;
  assign entries_vpn_p1__T_17_data = 10'h0;
  assign entries_vpn_p1__T_17_addr = 5'he;
  assign entries_vpn_p1__T_17_mask = 1'h0;
  assign entries_vpn_p1__T_17_en = reset | _T_1;
  assign entries_vpn_p1__T_18_data = 10'h0;
  assign entries_vpn_p1__T_18_addr = 5'hf;
  assign entries_vpn_p1__T_18_mask = 1'h0;
  assign entries_vpn_p1__T_18_en = reset | _T_1;
  assign entries_vpn_p1__T_19_data = 10'h0;
  assign entries_vpn_p1__T_19_addr = 5'h10;
  assign entries_vpn_p1__T_19_mask = 1'h0;
  assign entries_vpn_p1__T_19_en = reset | _T_1;
  assign entries_vpn_p1__T_20_data = 10'h0;
  assign entries_vpn_p1__T_20_addr = 5'h11;
  assign entries_vpn_p1__T_20_mask = 1'h0;
  assign entries_vpn_p1__T_20_en = reset | _T_1;
  assign entries_vpn_p1__T_21_data = 10'h0;
  assign entries_vpn_p1__T_21_addr = 5'h12;
  assign entries_vpn_p1__T_21_mask = 1'h0;
  assign entries_vpn_p1__T_21_en = reset | _T_1;
  assign entries_vpn_p1__T_22_data = 10'h0;
  assign entries_vpn_p1__T_22_addr = 5'h13;
  assign entries_vpn_p1__T_22_mask = 1'h0;
  assign entries_vpn_p1__T_22_en = reset | _T_1;
  assign entries_vpn_p1__T_23_data = 10'h0;
  assign entries_vpn_p1__T_23_addr = 5'h14;
  assign entries_vpn_p1__T_23_mask = 1'h0;
  assign entries_vpn_p1__T_23_en = reset | _T_1;
  assign entries_vpn_p1__T_24_data = 10'h0;
  assign entries_vpn_p1__T_24_addr = 5'h15;
  assign entries_vpn_p1__T_24_mask = 1'h0;
  assign entries_vpn_p1__T_24_en = reset | _T_1;
  assign entries_vpn_p1__T_25_data = 10'h0;
  assign entries_vpn_p1__T_25_addr = 5'h16;
  assign entries_vpn_p1__T_25_mask = 1'h0;
  assign entries_vpn_p1__T_25_en = reset | _T_1;
  assign entries_vpn_p1__T_26_data = 10'h0;
  assign entries_vpn_p1__T_26_addr = 5'h17;
  assign entries_vpn_p1__T_26_mask = 1'h0;
  assign entries_vpn_p1__T_26_en = reset | _T_1;
  assign entries_vpn_p1__T_27_data = 10'h0;
  assign entries_vpn_p1__T_27_addr = 5'h18;
  assign entries_vpn_p1__T_27_mask = 1'h0;
  assign entries_vpn_p1__T_27_en = reset | _T_1;
  assign entries_vpn_p1__T_28_data = 10'h0;
  assign entries_vpn_p1__T_28_addr = 5'h19;
  assign entries_vpn_p1__T_28_mask = 1'h0;
  assign entries_vpn_p1__T_28_en = reset | _T_1;
  assign entries_vpn_p1__T_29_data = 10'h0;
  assign entries_vpn_p1__T_29_addr = 5'h1a;
  assign entries_vpn_p1__T_29_mask = 1'h0;
  assign entries_vpn_p1__T_29_en = reset | _T_1;
  assign entries_vpn_p1__T_30_data = 10'h0;
  assign entries_vpn_p1__T_30_addr = 5'h1b;
  assign entries_vpn_p1__T_30_mask = 1'h0;
  assign entries_vpn_p1__T_30_en = reset | _T_1;
  assign entries_vpn_p1__T_31_data = 10'h0;
  assign entries_vpn_p1__T_31_addr = 5'h1c;
  assign entries_vpn_p1__T_31_mask = 1'h0;
  assign entries_vpn_p1__T_31_en = reset | _T_1;
  assign entries_vpn_p1__T_32_data = 10'h0;
  assign entries_vpn_p1__T_32_addr = 5'h1d;
  assign entries_vpn_p1__T_32_mask = 1'h0;
  assign entries_vpn_p1__T_32_en = reset | _T_1;
  assign entries_vpn_p1__T_33_data = 10'h0;
  assign entries_vpn_p1__T_33_addr = 5'h1e;
  assign entries_vpn_p1__T_33_mask = 1'h0;
  assign entries_vpn_p1__T_33_en = reset | _T_1;
  assign entries_vpn_p1__T_34_data = 10'h0;
  assign entries_vpn_p1__T_34_addr = 5'h1f;
  assign entries_vpn_p1__T_34_mask = 1'h0;
  assign entries_vpn_p1__T_34_en = reset | _T_1;
  assign entries_vpn_p1__T_57_data = 10'h0;
  assign entries_vpn_p1__T_57_addr = _T_55[4:0];
  assign entries_vpn_p1__T_57_mask = 1'h0;
  assign entries_vpn_p1__T_57_en = io_modify_mode == 2'h1;
  assign entries_vpn_p1__T_58_data = io_modify_vpn_p1;
  assign entries_vpn_p1__T_58_addr = _T_55[4:0];
  assign entries_vpn_p1__T_58_mask = 1'h1;
  assign entries_vpn_p1__T_58_en = io_modify_mode == 2'h1;
  assign entries_vpn_p1__T_59_data = 10'h0;
  assign entries_vpn_p1__T_59_addr = _T_55[4:0];
  assign entries_vpn_p1__T_59_mask = 1'h0;
  assign entries_vpn_p1__T_59_en = io_modify_mode == 2'h1;
  assign entries_vpn_p1__T_65_data = 10'h0;
  assign entries_vpn_p1__T_65_addr = _T_55[4:0];
  assign entries_vpn_p1__T_65_mask = 1'h0;
  assign entries_vpn_p1__T_65_en = _T_60 & _T_64;
  assign entries_pte_ppn_p2__T_39_addr = _T_37[4:0];
  assign entries_pte_ppn_p2__T_39_data = entries_pte_ppn_p2[entries_pte_ppn_p2__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p2__T_49_addr = _T_47[4:0];
  assign entries_pte_ppn_p2__T_49_data = entries_pte_ppn_p2[entries_pte_ppn_p2__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p2__T_61_addr = _T_55[4:0];
  assign entries_pte_ppn_p2__T_61_data = entries_pte_ppn_p2[entries_pte_ppn_p2__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p2__T_3_data = 10'h0;
  assign entries_pte_ppn_p2__T_3_addr = 5'h0;
  assign entries_pte_ppn_p2__T_3_mask = 1'h0;
  assign entries_pte_ppn_p2__T_3_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_4_data = 10'h0;
  assign entries_pte_ppn_p2__T_4_addr = 5'h1;
  assign entries_pte_ppn_p2__T_4_mask = 1'h0;
  assign entries_pte_ppn_p2__T_4_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_5_data = 10'h0;
  assign entries_pte_ppn_p2__T_5_addr = 5'h2;
  assign entries_pte_ppn_p2__T_5_mask = 1'h0;
  assign entries_pte_ppn_p2__T_5_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_6_data = 10'h0;
  assign entries_pte_ppn_p2__T_6_addr = 5'h3;
  assign entries_pte_ppn_p2__T_6_mask = 1'h0;
  assign entries_pte_ppn_p2__T_6_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_7_data = 10'h0;
  assign entries_pte_ppn_p2__T_7_addr = 5'h4;
  assign entries_pte_ppn_p2__T_7_mask = 1'h0;
  assign entries_pte_ppn_p2__T_7_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_8_data = 10'h0;
  assign entries_pte_ppn_p2__T_8_addr = 5'h5;
  assign entries_pte_ppn_p2__T_8_mask = 1'h0;
  assign entries_pte_ppn_p2__T_8_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_9_data = 10'h0;
  assign entries_pte_ppn_p2__T_9_addr = 5'h6;
  assign entries_pte_ppn_p2__T_9_mask = 1'h0;
  assign entries_pte_ppn_p2__T_9_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_10_data = 10'h0;
  assign entries_pte_ppn_p2__T_10_addr = 5'h7;
  assign entries_pte_ppn_p2__T_10_mask = 1'h0;
  assign entries_pte_ppn_p2__T_10_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_11_data = 10'h0;
  assign entries_pte_ppn_p2__T_11_addr = 5'h8;
  assign entries_pte_ppn_p2__T_11_mask = 1'h0;
  assign entries_pte_ppn_p2__T_11_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_12_data = 10'h0;
  assign entries_pte_ppn_p2__T_12_addr = 5'h9;
  assign entries_pte_ppn_p2__T_12_mask = 1'h0;
  assign entries_pte_ppn_p2__T_12_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_13_data = 10'h0;
  assign entries_pte_ppn_p2__T_13_addr = 5'ha;
  assign entries_pte_ppn_p2__T_13_mask = 1'h0;
  assign entries_pte_ppn_p2__T_13_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_14_data = 10'h0;
  assign entries_pte_ppn_p2__T_14_addr = 5'hb;
  assign entries_pte_ppn_p2__T_14_mask = 1'h0;
  assign entries_pte_ppn_p2__T_14_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_15_data = 10'h0;
  assign entries_pte_ppn_p2__T_15_addr = 5'hc;
  assign entries_pte_ppn_p2__T_15_mask = 1'h0;
  assign entries_pte_ppn_p2__T_15_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_16_data = 10'h0;
  assign entries_pte_ppn_p2__T_16_addr = 5'hd;
  assign entries_pte_ppn_p2__T_16_mask = 1'h0;
  assign entries_pte_ppn_p2__T_16_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_17_data = 10'h0;
  assign entries_pte_ppn_p2__T_17_addr = 5'he;
  assign entries_pte_ppn_p2__T_17_mask = 1'h0;
  assign entries_pte_ppn_p2__T_17_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_18_data = 10'h0;
  assign entries_pte_ppn_p2__T_18_addr = 5'hf;
  assign entries_pte_ppn_p2__T_18_mask = 1'h0;
  assign entries_pte_ppn_p2__T_18_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_19_data = 10'h0;
  assign entries_pte_ppn_p2__T_19_addr = 5'h10;
  assign entries_pte_ppn_p2__T_19_mask = 1'h0;
  assign entries_pte_ppn_p2__T_19_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_20_data = 10'h0;
  assign entries_pte_ppn_p2__T_20_addr = 5'h11;
  assign entries_pte_ppn_p2__T_20_mask = 1'h0;
  assign entries_pte_ppn_p2__T_20_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_21_data = 10'h0;
  assign entries_pte_ppn_p2__T_21_addr = 5'h12;
  assign entries_pte_ppn_p2__T_21_mask = 1'h0;
  assign entries_pte_ppn_p2__T_21_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_22_data = 10'h0;
  assign entries_pte_ppn_p2__T_22_addr = 5'h13;
  assign entries_pte_ppn_p2__T_22_mask = 1'h0;
  assign entries_pte_ppn_p2__T_22_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_23_data = 10'h0;
  assign entries_pte_ppn_p2__T_23_addr = 5'h14;
  assign entries_pte_ppn_p2__T_23_mask = 1'h0;
  assign entries_pte_ppn_p2__T_23_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_24_data = 10'h0;
  assign entries_pte_ppn_p2__T_24_addr = 5'h15;
  assign entries_pte_ppn_p2__T_24_mask = 1'h0;
  assign entries_pte_ppn_p2__T_24_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_25_data = 10'h0;
  assign entries_pte_ppn_p2__T_25_addr = 5'h16;
  assign entries_pte_ppn_p2__T_25_mask = 1'h0;
  assign entries_pte_ppn_p2__T_25_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_26_data = 10'h0;
  assign entries_pte_ppn_p2__T_26_addr = 5'h17;
  assign entries_pte_ppn_p2__T_26_mask = 1'h0;
  assign entries_pte_ppn_p2__T_26_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_27_data = 10'h0;
  assign entries_pte_ppn_p2__T_27_addr = 5'h18;
  assign entries_pte_ppn_p2__T_27_mask = 1'h0;
  assign entries_pte_ppn_p2__T_27_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_28_data = 10'h0;
  assign entries_pte_ppn_p2__T_28_addr = 5'h19;
  assign entries_pte_ppn_p2__T_28_mask = 1'h0;
  assign entries_pte_ppn_p2__T_28_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_29_data = 10'h0;
  assign entries_pte_ppn_p2__T_29_addr = 5'h1a;
  assign entries_pte_ppn_p2__T_29_mask = 1'h0;
  assign entries_pte_ppn_p2__T_29_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_30_data = 10'h0;
  assign entries_pte_ppn_p2__T_30_addr = 5'h1b;
  assign entries_pte_ppn_p2__T_30_mask = 1'h0;
  assign entries_pte_ppn_p2__T_30_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_31_data = 10'h0;
  assign entries_pte_ppn_p2__T_31_addr = 5'h1c;
  assign entries_pte_ppn_p2__T_31_mask = 1'h0;
  assign entries_pte_ppn_p2__T_31_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_32_data = 10'h0;
  assign entries_pte_ppn_p2__T_32_addr = 5'h1d;
  assign entries_pte_ppn_p2__T_32_mask = 1'h0;
  assign entries_pte_ppn_p2__T_32_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_33_data = 10'h0;
  assign entries_pte_ppn_p2__T_33_addr = 5'h1e;
  assign entries_pte_ppn_p2__T_33_mask = 1'h0;
  assign entries_pte_ppn_p2__T_33_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_34_data = 10'h0;
  assign entries_pte_ppn_p2__T_34_addr = 5'h1f;
  assign entries_pte_ppn_p2__T_34_mask = 1'h0;
  assign entries_pte_ppn_p2__T_34_en = reset | _T_1;
  assign entries_pte_ppn_p2__T_57_data = 10'h0;
  assign entries_pte_ppn_p2__T_57_addr = _T_55[4:0];
  assign entries_pte_ppn_p2__T_57_mask = 1'h0;
  assign entries_pte_ppn_p2__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p2__T_58_data = 10'h0;
  assign entries_pte_ppn_p2__T_58_addr = _T_55[4:0];
  assign entries_pte_ppn_p2__T_58_mask = 1'h0;
  assign entries_pte_ppn_p2__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p2__T_59_data = io_modify_pte_ppn_p2;
  assign entries_pte_ppn_p2__T_59_addr = _T_55[4:0];
  assign entries_pte_ppn_p2__T_59_mask = 1'h1;
  assign entries_pte_ppn_p2__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p2__T_65_data = 10'h0;
  assign entries_pte_ppn_p2__T_65_addr = _T_55[4:0];
  assign entries_pte_ppn_p2__T_65_mask = 1'h0;
  assign entries_pte_ppn_p2__T_65_en = _T_60 & _T_64;
  assign entries_pte_ppn_p1__T_39_addr = _T_37[4:0];
  assign entries_pte_ppn_p1__T_39_data = entries_pte_ppn_p1[entries_pte_ppn_p1__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p1__T_49_addr = _T_47[4:0];
  assign entries_pte_ppn_p1__T_49_data = entries_pte_ppn_p1[entries_pte_ppn_p1__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p1__T_61_addr = _T_55[4:0];
  assign entries_pte_ppn_p1__T_61_data = entries_pte_ppn_p1[entries_pte_ppn_p1__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_ppn_p1__T_3_data = 10'h0;
  assign entries_pte_ppn_p1__T_3_addr = 5'h0;
  assign entries_pte_ppn_p1__T_3_mask = 1'h0;
  assign entries_pte_ppn_p1__T_3_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_4_data = 10'h0;
  assign entries_pte_ppn_p1__T_4_addr = 5'h1;
  assign entries_pte_ppn_p1__T_4_mask = 1'h0;
  assign entries_pte_ppn_p1__T_4_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_5_data = 10'h0;
  assign entries_pte_ppn_p1__T_5_addr = 5'h2;
  assign entries_pte_ppn_p1__T_5_mask = 1'h0;
  assign entries_pte_ppn_p1__T_5_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_6_data = 10'h0;
  assign entries_pte_ppn_p1__T_6_addr = 5'h3;
  assign entries_pte_ppn_p1__T_6_mask = 1'h0;
  assign entries_pte_ppn_p1__T_6_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_7_data = 10'h0;
  assign entries_pte_ppn_p1__T_7_addr = 5'h4;
  assign entries_pte_ppn_p1__T_7_mask = 1'h0;
  assign entries_pte_ppn_p1__T_7_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_8_data = 10'h0;
  assign entries_pte_ppn_p1__T_8_addr = 5'h5;
  assign entries_pte_ppn_p1__T_8_mask = 1'h0;
  assign entries_pte_ppn_p1__T_8_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_9_data = 10'h0;
  assign entries_pte_ppn_p1__T_9_addr = 5'h6;
  assign entries_pte_ppn_p1__T_9_mask = 1'h0;
  assign entries_pte_ppn_p1__T_9_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_10_data = 10'h0;
  assign entries_pte_ppn_p1__T_10_addr = 5'h7;
  assign entries_pte_ppn_p1__T_10_mask = 1'h0;
  assign entries_pte_ppn_p1__T_10_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_11_data = 10'h0;
  assign entries_pte_ppn_p1__T_11_addr = 5'h8;
  assign entries_pte_ppn_p1__T_11_mask = 1'h0;
  assign entries_pte_ppn_p1__T_11_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_12_data = 10'h0;
  assign entries_pte_ppn_p1__T_12_addr = 5'h9;
  assign entries_pte_ppn_p1__T_12_mask = 1'h0;
  assign entries_pte_ppn_p1__T_12_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_13_data = 10'h0;
  assign entries_pte_ppn_p1__T_13_addr = 5'ha;
  assign entries_pte_ppn_p1__T_13_mask = 1'h0;
  assign entries_pte_ppn_p1__T_13_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_14_data = 10'h0;
  assign entries_pte_ppn_p1__T_14_addr = 5'hb;
  assign entries_pte_ppn_p1__T_14_mask = 1'h0;
  assign entries_pte_ppn_p1__T_14_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_15_data = 10'h0;
  assign entries_pte_ppn_p1__T_15_addr = 5'hc;
  assign entries_pte_ppn_p1__T_15_mask = 1'h0;
  assign entries_pte_ppn_p1__T_15_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_16_data = 10'h0;
  assign entries_pte_ppn_p1__T_16_addr = 5'hd;
  assign entries_pte_ppn_p1__T_16_mask = 1'h0;
  assign entries_pte_ppn_p1__T_16_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_17_data = 10'h0;
  assign entries_pte_ppn_p1__T_17_addr = 5'he;
  assign entries_pte_ppn_p1__T_17_mask = 1'h0;
  assign entries_pte_ppn_p1__T_17_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_18_data = 10'h0;
  assign entries_pte_ppn_p1__T_18_addr = 5'hf;
  assign entries_pte_ppn_p1__T_18_mask = 1'h0;
  assign entries_pte_ppn_p1__T_18_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_19_data = 10'h0;
  assign entries_pte_ppn_p1__T_19_addr = 5'h10;
  assign entries_pte_ppn_p1__T_19_mask = 1'h0;
  assign entries_pte_ppn_p1__T_19_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_20_data = 10'h0;
  assign entries_pte_ppn_p1__T_20_addr = 5'h11;
  assign entries_pte_ppn_p1__T_20_mask = 1'h0;
  assign entries_pte_ppn_p1__T_20_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_21_data = 10'h0;
  assign entries_pte_ppn_p1__T_21_addr = 5'h12;
  assign entries_pte_ppn_p1__T_21_mask = 1'h0;
  assign entries_pte_ppn_p1__T_21_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_22_data = 10'h0;
  assign entries_pte_ppn_p1__T_22_addr = 5'h13;
  assign entries_pte_ppn_p1__T_22_mask = 1'h0;
  assign entries_pte_ppn_p1__T_22_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_23_data = 10'h0;
  assign entries_pte_ppn_p1__T_23_addr = 5'h14;
  assign entries_pte_ppn_p1__T_23_mask = 1'h0;
  assign entries_pte_ppn_p1__T_23_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_24_data = 10'h0;
  assign entries_pte_ppn_p1__T_24_addr = 5'h15;
  assign entries_pte_ppn_p1__T_24_mask = 1'h0;
  assign entries_pte_ppn_p1__T_24_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_25_data = 10'h0;
  assign entries_pte_ppn_p1__T_25_addr = 5'h16;
  assign entries_pte_ppn_p1__T_25_mask = 1'h0;
  assign entries_pte_ppn_p1__T_25_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_26_data = 10'h0;
  assign entries_pte_ppn_p1__T_26_addr = 5'h17;
  assign entries_pte_ppn_p1__T_26_mask = 1'h0;
  assign entries_pte_ppn_p1__T_26_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_27_data = 10'h0;
  assign entries_pte_ppn_p1__T_27_addr = 5'h18;
  assign entries_pte_ppn_p1__T_27_mask = 1'h0;
  assign entries_pte_ppn_p1__T_27_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_28_data = 10'h0;
  assign entries_pte_ppn_p1__T_28_addr = 5'h19;
  assign entries_pte_ppn_p1__T_28_mask = 1'h0;
  assign entries_pte_ppn_p1__T_28_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_29_data = 10'h0;
  assign entries_pte_ppn_p1__T_29_addr = 5'h1a;
  assign entries_pte_ppn_p1__T_29_mask = 1'h0;
  assign entries_pte_ppn_p1__T_29_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_30_data = 10'h0;
  assign entries_pte_ppn_p1__T_30_addr = 5'h1b;
  assign entries_pte_ppn_p1__T_30_mask = 1'h0;
  assign entries_pte_ppn_p1__T_30_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_31_data = 10'h0;
  assign entries_pte_ppn_p1__T_31_addr = 5'h1c;
  assign entries_pte_ppn_p1__T_31_mask = 1'h0;
  assign entries_pte_ppn_p1__T_31_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_32_data = 10'h0;
  assign entries_pte_ppn_p1__T_32_addr = 5'h1d;
  assign entries_pte_ppn_p1__T_32_mask = 1'h0;
  assign entries_pte_ppn_p1__T_32_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_33_data = 10'h0;
  assign entries_pte_ppn_p1__T_33_addr = 5'h1e;
  assign entries_pte_ppn_p1__T_33_mask = 1'h0;
  assign entries_pte_ppn_p1__T_33_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_34_data = 10'h0;
  assign entries_pte_ppn_p1__T_34_addr = 5'h1f;
  assign entries_pte_ppn_p1__T_34_mask = 1'h0;
  assign entries_pte_ppn_p1__T_34_en = reset | _T_1;
  assign entries_pte_ppn_p1__T_57_data = 10'h0;
  assign entries_pte_ppn_p1__T_57_addr = _T_55[4:0];
  assign entries_pte_ppn_p1__T_57_mask = 1'h0;
  assign entries_pte_ppn_p1__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p1__T_58_data = 10'h0;
  assign entries_pte_ppn_p1__T_58_addr = _T_55[4:0];
  assign entries_pte_ppn_p1__T_58_mask = 1'h0;
  assign entries_pte_ppn_p1__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p1__T_59_data = io_modify_pte_ppn_p1;
  assign entries_pte_ppn_p1__T_59_addr = _T_55[4:0];
  assign entries_pte_ppn_p1__T_59_mask = 1'h1;
  assign entries_pte_ppn_p1__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_ppn_p1__T_65_data = 10'h0;
  assign entries_pte_ppn_p1__T_65_addr = _T_55[4:0];
  assign entries_pte_ppn_p1__T_65_mask = 1'h0;
  assign entries_pte_ppn_p1__T_65_en = _T_60 & _T_64;
  assign entries_pte_U__T_39_addr = _T_37[4:0];
  assign entries_pte_U__T_39_data = entries_pte_U[entries_pte_U__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_U__T_49_addr = _T_47[4:0];
  assign entries_pte_U__T_49_data = entries_pte_U[entries_pte_U__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_U__T_61_addr = _T_55[4:0];
  assign entries_pte_U__T_61_data = entries_pte_U[entries_pte_U__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_U__T_3_data = 1'h0;
  assign entries_pte_U__T_3_addr = 5'h0;
  assign entries_pte_U__T_3_mask = 1'h0;
  assign entries_pte_U__T_3_en = reset | _T_1;
  assign entries_pte_U__T_4_data = 1'h0;
  assign entries_pte_U__T_4_addr = 5'h1;
  assign entries_pte_U__T_4_mask = 1'h0;
  assign entries_pte_U__T_4_en = reset | _T_1;
  assign entries_pte_U__T_5_data = 1'h0;
  assign entries_pte_U__T_5_addr = 5'h2;
  assign entries_pte_U__T_5_mask = 1'h0;
  assign entries_pte_U__T_5_en = reset | _T_1;
  assign entries_pte_U__T_6_data = 1'h0;
  assign entries_pte_U__T_6_addr = 5'h3;
  assign entries_pte_U__T_6_mask = 1'h0;
  assign entries_pte_U__T_6_en = reset | _T_1;
  assign entries_pte_U__T_7_data = 1'h0;
  assign entries_pte_U__T_7_addr = 5'h4;
  assign entries_pte_U__T_7_mask = 1'h0;
  assign entries_pte_U__T_7_en = reset | _T_1;
  assign entries_pte_U__T_8_data = 1'h0;
  assign entries_pte_U__T_8_addr = 5'h5;
  assign entries_pte_U__T_8_mask = 1'h0;
  assign entries_pte_U__T_8_en = reset | _T_1;
  assign entries_pte_U__T_9_data = 1'h0;
  assign entries_pte_U__T_9_addr = 5'h6;
  assign entries_pte_U__T_9_mask = 1'h0;
  assign entries_pte_U__T_9_en = reset | _T_1;
  assign entries_pte_U__T_10_data = 1'h0;
  assign entries_pte_U__T_10_addr = 5'h7;
  assign entries_pte_U__T_10_mask = 1'h0;
  assign entries_pte_U__T_10_en = reset | _T_1;
  assign entries_pte_U__T_11_data = 1'h0;
  assign entries_pte_U__T_11_addr = 5'h8;
  assign entries_pte_U__T_11_mask = 1'h0;
  assign entries_pte_U__T_11_en = reset | _T_1;
  assign entries_pte_U__T_12_data = 1'h0;
  assign entries_pte_U__T_12_addr = 5'h9;
  assign entries_pte_U__T_12_mask = 1'h0;
  assign entries_pte_U__T_12_en = reset | _T_1;
  assign entries_pte_U__T_13_data = 1'h0;
  assign entries_pte_U__T_13_addr = 5'ha;
  assign entries_pte_U__T_13_mask = 1'h0;
  assign entries_pte_U__T_13_en = reset | _T_1;
  assign entries_pte_U__T_14_data = 1'h0;
  assign entries_pte_U__T_14_addr = 5'hb;
  assign entries_pte_U__T_14_mask = 1'h0;
  assign entries_pte_U__T_14_en = reset | _T_1;
  assign entries_pte_U__T_15_data = 1'h0;
  assign entries_pte_U__T_15_addr = 5'hc;
  assign entries_pte_U__T_15_mask = 1'h0;
  assign entries_pte_U__T_15_en = reset | _T_1;
  assign entries_pte_U__T_16_data = 1'h0;
  assign entries_pte_U__T_16_addr = 5'hd;
  assign entries_pte_U__T_16_mask = 1'h0;
  assign entries_pte_U__T_16_en = reset | _T_1;
  assign entries_pte_U__T_17_data = 1'h0;
  assign entries_pte_U__T_17_addr = 5'he;
  assign entries_pte_U__T_17_mask = 1'h0;
  assign entries_pte_U__T_17_en = reset | _T_1;
  assign entries_pte_U__T_18_data = 1'h0;
  assign entries_pte_U__T_18_addr = 5'hf;
  assign entries_pte_U__T_18_mask = 1'h0;
  assign entries_pte_U__T_18_en = reset | _T_1;
  assign entries_pte_U__T_19_data = 1'h0;
  assign entries_pte_U__T_19_addr = 5'h10;
  assign entries_pte_U__T_19_mask = 1'h0;
  assign entries_pte_U__T_19_en = reset | _T_1;
  assign entries_pte_U__T_20_data = 1'h0;
  assign entries_pte_U__T_20_addr = 5'h11;
  assign entries_pte_U__T_20_mask = 1'h0;
  assign entries_pte_U__T_20_en = reset | _T_1;
  assign entries_pte_U__T_21_data = 1'h0;
  assign entries_pte_U__T_21_addr = 5'h12;
  assign entries_pte_U__T_21_mask = 1'h0;
  assign entries_pte_U__T_21_en = reset | _T_1;
  assign entries_pte_U__T_22_data = 1'h0;
  assign entries_pte_U__T_22_addr = 5'h13;
  assign entries_pte_U__T_22_mask = 1'h0;
  assign entries_pte_U__T_22_en = reset | _T_1;
  assign entries_pte_U__T_23_data = 1'h0;
  assign entries_pte_U__T_23_addr = 5'h14;
  assign entries_pte_U__T_23_mask = 1'h0;
  assign entries_pte_U__T_23_en = reset | _T_1;
  assign entries_pte_U__T_24_data = 1'h0;
  assign entries_pte_U__T_24_addr = 5'h15;
  assign entries_pte_U__T_24_mask = 1'h0;
  assign entries_pte_U__T_24_en = reset | _T_1;
  assign entries_pte_U__T_25_data = 1'h0;
  assign entries_pte_U__T_25_addr = 5'h16;
  assign entries_pte_U__T_25_mask = 1'h0;
  assign entries_pte_U__T_25_en = reset | _T_1;
  assign entries_pte_U__T_26_data = 1'h0;
  assign entries_pte_U__T_26_addr = 5'h17;
  assign entries_pte_U__T_26_mask = 1'h0;
  assign entries_pte_U__T_26_en = reset | _T_1;
  assign entries_pte_U__T_27_data = 1'h0;
  assign entries_pte_U__T_27_addr = 5'h18;
  assign entries_pte_U__T_27_mask = 1'h0;
  assign entries_pte_U__T_27_en = reset | _T_1;
  assign entries_pte_U__T_28_data = 1'h0;
  assign entries_pte_U__T_28_addr = 5'h19;
  assign entries_pte_U__T_28_mask = 1'h0;
  assign entries_pte_U__T_28_en = reset | _T_1;
  assign entries_pte_U__T_29_data = 1'h0;
  assign entries_pte_U__T_29_addr = 5'h1a;
  assign entries_pte_U__T_29_mask = 1'h0;
  assign entries_pte_U__T_29_en = reset | _T_1;
  assign entries_pte_U__T_30_data = 1'h0;
  assign entries_pte_U__T_30_addr = 5'h1b;
  assign entries_pte_U__T_30_mask = 1'h0;
  assign entries_pte_U__T_30_en = reset | _T_1;
  assign entries_pte_U__T_31_data = 1'h0;
  assign entries_pte_U__T_31_addr = 5'h1c;
  assign entries_pte_U__T_31_mask = 1'h0;
  assign entries_pte_U__T_31_en = reset | _T_1;
  assign entries_pte_U__T_32_data = 1'h0;
  assign entries_pte_U__T_32_addr = 5'h1d;
  assign entries_pte_U__T_32_mask = 1'h0;
  assign entries_pte_U__T_32_en = reset | _T_1;
  assign entries_pte_U__T_33_data = 1'h0;
  assign entries_pte_U__T_33_addr = 5'h1e;
  assign entries_pte_U__T_33_mask = 1'h0;
  assign entries_pte_U__T_33_en = reset | _T_1;
  assign entries_pte_U__T_34_data = 1'h0;
  assign entries_pte_U__T_34_addr = 5'h1f;
  assign entries_pte_U__T_34_mask = 1'h0;
  assign entries_pte_U__T_34_en = reset | _T_1;
  assign entries_pte_U__T_57_data = 1'h0;
  assign entries_pte_U__T_57_addr = _T_55[4:0];
  assign entries_pte_U__T_57_mask = 1'h0;
  assign entries_pte_U__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_U__T_58_data = 1'h0;
  assign entries_pte_U__T_58_addr = _T_55[4:0];
  assign entries_pte_U__T_58_mask = 1'h0;
  assign entries_pte_U__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_U__T_59_data = io_modify_pte_U;
  assign entries_pte_U__T_59_addr = _T_55[4:0];
  assign entries_pte_U__T_59_mask = 1'h1;
  assign entries_pte_U__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_U__T_65_data = 1'h0;
  assign entries_pte_U__T_65_addr = _T_55[4:0];
  assign entries_pte_U__T_65_mask = 1'h0;
  assign entries_pte_U__T_65_en = _T_60 & _T_64;
  assign entries_pte_X__T_39_addr = _T_37[4:0];
  assign entries_pte_X__T_39_data = entries_pte_X[entries_pte_X__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_X__T_49_addr = _T_47[4:0];
  assign entries_pte_X__T_49_data = entries_pte_X[entries_pte_X__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_X__T_61_addr = _T_55[4:0];
  assign entries_pte_X__T_61_data = entries_pte_X[entries_pte_X__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_X__T_3_data = 1'h0;
  assign entries_pte_X__T_3_addr = 5'h0;
  assign entries_pte_X__T_3_mask = 1'h0;
  assign entries_pte_X__T_3_en = reset | _T_1;
  assign entries_pte_X__T_4_data = 1'h0;
  assign entries_pte_X__T_4_addr = 5'h1;
  assign entries_pte_X__T_4_mask = 1'h0;
  assign entries_pte_X__T_4_en = reset | _T_1;
  assign entries_pte_X__T_5_data = 1'h0;
  assign entries_pte_X__T_5_addr = 5'h2;
  assign entries_pte_X__T_5_mask = 1'h0;
  assign entries_pte_X__T_5_en = reset | _T_1;
  assign entries_pte_X__T_6_data = 1'h0;
  assign entries_pte_X__T_6_addr = 5'h3;
  assign entries_pte_X__T_6_mask = 1'h0;
  assign entries_pte_X__T_6_en = reset | _T_1;
  assign entries_pte_X__T_7_data = 1'h0;
  assign entries_pte_X__T_7_addr = 5'h4;
  assign entries_pte_X__T_7_mask = 1'h0;
  assign entries_pte_X__T_7_en = reset | _T_1;
  assign entries_pte_X__T_8_data = 1'h0;
  assign entries_pte_X__T_8_addr = 5'h5;
  assign entries_pte_X__T_8_mask = 1'h0;
  assign entries_pte_X__T_8_en = reset | _T_1;
  assign entries_pte_X__T_9_data = 1'h0;
  assign entries_pte_X__T_9_addr = 5'h6;
  assign entries_pte_X__T_9_mask = 1'h0;
  assign entries_pte_X__T_9_en = reset | _T_1;
  assign entries_pte_X__T_10_data = 1'h0;
  assign entries_pte_X__T_10_addr = 5'h7;
  assign entries_pte_X__T_10_mask = 1'h0;
  assign entries_pte_X__T_10_en = reset | _T_1;
  assign entries_pte_X__T_11_data = 1'h0;
  assign entries_pte_X__T_11_addr = 5'h8;
  assign entries_pte_X__T_11_mask = 1'h0;
  assign entries_pte_X__T_11_en = reset | _T_1;
  assign entries_pte_X__T_12_data = 1'h0;
  assign entries_pte_X__T_12_addr = 5'h9;
  assign entries_pte_X__T_12_mask = 1'h0;
  assign entries_pte_X__T_12_en = reset | _T_1;
  assign entries_pte_X__T_13_data = 1'h0;
  assign entries_pte_X__T_13_addr = 5'ha;
  assign entries_pte_X__T_13_mask = 1'h0;
  assign entries_pte_X__T_13_en = reset | _T_1;
  assign entries_pte_X__T_14_data = 1'h0;
  assign entries_pte_X__T_14_addr = 5'hb;
  assign entries_pte_X__T_14_mask = 1'h0;
  assign entries_pte_X__T_14_en = reset | _T_1;
  assign entries_pte_X__T_15_data = 1'h0;
  assign entries_pte_X__T_15_addr = 5'hc;
  assign entries_pte_X__T_15_mask = 1'h0;
  assign entries_pte_X__T_15_en = reset | _T_1;
  assign entries_pte_X__T_16_data = 1'h0;
  assign entries_pte_X__T_16_addr = 5'hd;
  assign entries_pte_X__T_16_mask = 1'h0;
  assign entries_pte_X__T_16_en = reset | _T_1;
  assign entries_pte_X__T_17_data = 1'h0;
  assign entries_pte_X__T_17_addr = 5'he;
  assign entries_pte_X__T_17_mask = 1'h0;
  assign entries_pte_X__T_17_en = reset | _T_1;
  assign entries_pte_X__T_18_data = 1'h0;
  assign entries_pte_X__T_18_addr = 5'hf;
  assign entries_pte_X__T_18_mask = 1'h0;
  assign entries_pte_X__T_18_en = reset | _T_1;
  assign entries_pte_X__T_19_data = 1'h0;
  assign entries_pte_X__T_19_addr = 5'h10;
  assign entries_pte_X__T_19_mask = 1'h0;
  assign entries_pte_X__T_19_en = reset | _T_1;
  assign entries_pte_X__T_20_data = 1'h0;
  assign entries_pte_X__T_20_addr = 5'h11;
  assign entries_pte_X__T_20_mask = 1'h0;
  assign entries_pte_X__T_20_en = reset | _T_1;
  assign entries_pte_X__T_21_data = 1'h0;
  assign entries_pte_X__T_21_addr = 5'h12;
  assign entries_pte_X__T_21_mask = 1'h0;
  assign entries_pte_X__T_21_en = reset | _T_1;
  assign entries_pte_X__T_22_data = 1'h0;
  assign entries_pte_X__T_22_addr = 5'h13;
  assign entries_pte_X__T_22_mask = 1'h0;
  assign entries_pte_X__T_22_en = reset | _T_1;
  assign entries_pte_X__T_23_data = 1'h0;
  assign entries_pte_X__T_23_addr = 5'h14;
  assign entries_pte_X__T_23_mask = 1'h0;
  assign entries_pte_X__T_23_en = reset | _T_1;
  assign entries_pte_X__T_24_data = 1'h0;
  assign entries_pte_X__T_24_addr = 5'h15;
  assign entries_pte_X__T_24_mask = 1'h0;
  assign entries_pte_X__T_24_en = reset | _T_1;
  assign entries_pte_X__T_25_data = 1'h0;
  assign entries_pte_X__T_25_addr = 5'h16;
  assign entries_pte_X__T_25_mask = 1'h0;
  assign entries_pte_X__T_25_en = reset | _T_1;
  assign entries_pte_X__T_26_data = 1'h0;
  assign entries_pte_X__T_26_addr = 5'h17;
  assign entries_pte_X__T_26_mask = 1'h0;
  assign entries_pte_X__T_26_en = reset | _T_1;
  assign entries_pte_X__T_27_data = 1'h0;
  assign entries_pte_X__T_27_addr = 5'h18;
  assign entries_pte_X__T_27_mask = 1'h0;
  assign entries_pte_X__T_27_en = reset | _T_1;
  assign entries_pte_X__T_28_data = 1'h0;
  assign entries_pte_X__T_28_addr = 5'h19;
  assign entries_pte_X__T_28_mask = 1'h0;
  assign entries_pte_X__T_28_en = reset | _T_1;
  assign entries_pte_X__T_29_data = 1'h0;
  assign entries_pte_X__T_29_addr = 5'h1a;
  assign entries_pte_X__T_29_mask = 1'h0;
  assign entries_pte_X__T_29_en = reset | _T_1;
  assign entries_pte_X__T_30_data = 1'h0;
  assign entries_pte_X__T_30_addr = 5'h1b;
  assign entries_pte_X__T_30_mask = 1'h0;
  assign entries_pte_X__T_30_en = reset | _T_1;
  assign entries_pte_X__T_31_data = 1'h0;
  assign entries_pte_X__T_31_addr = 5'h1c;
  assign entries_pte_X__T_31_mask = 1'h0;
  assign entries_pte_X__T_31_en = reset | _T_1;
  assign entries_pte_X__T_32_data = 1'h0;
  assign entries_pte_X__T_32_addr = 5'h1d;
  assign entries_pte_X__T_32_mask = 1'h0;
  assign entries_pte_X__T_32_en = reset | _T_1;
  assign entries_pte_X__T_33_data = 1'h0;
  assign entries_pte_X__T_33_addr = 5'h1e;
  assign entries_pte_X__T_33_mask = 1'h0;
  assign entries_pte_X__T_33_en = reset | _T_1;
  assign entries_pte_X__T_34_data = 1'h0;
  assign entries_pte_X__T_34_addr = 5'h1f;
  assign entries_pte_X__T_34_mask = 1'h0;
  assign entries_pte_X__T_34_en = reset | _T_1;
  assign entries_pte_X__T_57_data = 1'h0;
  assign entries_pte_X__T_57_addr = _T_55[4:0];
  assign entries_pte_X__T_57_mask = 1'h0;
  assign entries_pte_X__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_X__T_58_data = 1'h0;
  assign entries_pte_X__T_58_addr = _T_55[4:0];
  assign entries_pte_X__T_58_mask = 1'h0;
  assign entries_pte_X__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_X__T_59_data = io_modify_pte_X;
  assign entries_pte_X__T_59_addr = _T_55[4:0];
  assign entries_pte_X__T_59_mask = 1'h1;
  assign entries_pte_X__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_X__T_65_data = 1'h0;
  assign entries_pte_X__T_65_addr = _T_55[4:0];
  assign entries_pte_X__T_65_mask = 1'h0;
  assign entries_pte_X__T_65_en = _T_60 & _T_64;
  assign entries_pte_W__T_39_addr = _T_37[4:0];
  assign entries_pte_W__T_39_data = entries_pte_W[entries_pte_W__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_W__T_49_addr = _T_47[4:0];
  assign entries_pte_W__T_49_data = entries_pte_W[entries_pte_W__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_W__T_61_addr = _T_55[4:0];
  assign entries_pte_W__T_61_data = entries_pte_W[entries_pte_W__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_W__T_3_data = 1'h0;
  assign entries_pte_W__T_3_addr = 5'h0;
  assign entries_pte_W__T_3_mask = 1'h0;
  assign entries_pte_W__T_3_en = reset | _T_1;
  assign entries_pte_W__T_4_data = 1'h0;
  assign entries_pte_W__T_4_addr = 5'h1;
  assign entries_pte_W__T_4_mask = 1'h0;
  assign entries_pte_W__T_4_en = reset | _T_1;
  assign entries_pte_W__T_5_data = 1'h0;
  assign entries_pte_W__T_5_addr = 5'h2;
  assign entries_pte_W__T_5_mask = 1'h0;
  assign entries_pte_W__T_5_en = reset | _T_1;
  assign entries_pte_W__T_6_data = 1'h0;
  assign entries_pte_W__T_6_addr = 5'h3;
  assign entries_pte_W__T_6_mask = 1'h0;
  assign entries_pte_W__T_6_en = reset | _T_1;
  assign entries_pte_W__T_7_data = 1'h0;
  assign entries_pte_W__T_7_addr = 5'h4;
  assign entries_pte_W__T_7_mask = 1'h0;
  assign entries_pte_W__T_7_en = reset | _T_1;
  assign entries_pte_W__T_8_data = 1'h0;
  assign entries_pte_W__T_8_addr = 5'h5;
  assign entries_pte_W__T_8_mask = 1'h0;
  assign entries_pte_W__T_8_en = reset | _T_1;
  assign entries_pte_W__T_9_data = 1'h0;
  assign entries_pte_W__T_9_addr = 5'h6;
  assign entries_pte_W__T_9_mask = 1'h0;
  assign entries_pte_W__T_9_en = reset | _T_1;
  assign entries_pte_W__T_10_data = 1'h0;
  assign entries_pte_W__T_10_addr = 5'h7;
  assign entries_pte_W__T_10_mask = 1'h0;
  assign entries_pte_W__T_10_en = reset | _T_1;
  assign entries_pte_W__T_11_data = 1'h0;
  assign entries_pte_W__T_11_addr = 5'h8;
  assign entries_pte_W__T_11_mask = 1'h0;
  assign entries_pte_W__T_11_en = reset | _T_1;
  assign entries_pte_W__T_12_data = 1'h0;
  assign entries_pte_W__T_12_addr = 5'h9;
  assign entries_pte_W__T_12_mask = 1'h0;
  assign entries_pte_W__T_12_en = reset | _T_1;
  assign entries_pte_W__T_13_data = 1'h0;
  assign entries_pte_W__T_13_addr = 5'ha;
  assign entries_pte_W__T_13_mask = 1'h0;
  assign entries_pte_W__T_13_en = reset | _T_1;
  assign entries_pte_W__T_14_data = 1'h0;
  assign entries_pte_W__T_14_addr = 5'hb;
  assign entries_pte_W__T_14_mask = 1'h0;
  assign entries_pte_W__T_14_en = reset | _T_1;
  assign entries_pte_W__T_15_data = 1'h0;
  assign entries_pte_W__T_15_addr = 5'hc;
  assign entries_pte_W__T_15_mask = 1'h0;
  assign entries_pte_W__T_15_en = reset | _T_1;
  assign entries_pte_W__T_16_data = 1'h0;
  assign entries_pte_W__T_16_addr = 5'hd;
  assign entries_pte_W__T_16_mask = 1'h0;
  assign entries_pte_W__T_16_en = reset | _T_1;
  assign entries_pte_W__T_17_data = 1'h0;
  assign entries_pte_W__T_17_addr = 5'he;
  assign entries_pte_W__T_17_mask = 1'h0;
  assign entries_pte_W__T_17_en = reset | _T_1;
  assign entries_pte_W__T_18_data = 1'h0;
  assign entries_pte_W__T_18_addr = 5'hf;
  assign entries_pte_W__T_18_mask = 1'h0;
  assign entries_pte_W__T_18_en = reset | _T_1;
  assign entries_pte_W__T_19_data = 1'h0;
  assign entries_pte_W__T_19_addr = 5'h10;
  assign entries_pte_W__T_19_mask = 1'h0;
  assign entries_pte_W__T_19_en = reset | _T_1;
  assign entries_pte_W__T_20_data = 1'h0;
  assign entries_pte_W__T_20_addr = 5'h11;
  assign entries_pte_W__T_20_mask = 1'h0;
  assign entries_pte_W__T_20_en = reset | _T_1;
  assign entries_pte_W__T_21_data = 1'h0;
  assign entries_pte_W__T_21_addr = 5'h12;
  assign entries_pte_W__T_21_mask = 1'h0;
  assign entries_pte_W__T_21_en = reset | _T_1;
  assign entries_pte_W__T_22_data = 1'h0;
  assign entries_pte_W__T_22_addr = 5'h13;
  assign entries_pte_W__T_22_mask = 1'h0;
  assign entries_pte_W__T_22_en = reset | _T_1;
  assign entries_pte_W__T_23_data = 1'h0;
  assign entries_pte_W__T_23_addr = 5'h14;
  assign entries_pte_W__T_23_mask = 1'h0;
  assign entries_pte_W__T_23_en = reset | _T_1;
  assign entries_pte_W__T_24_data = 1'h0;
  assign entries_pte_W__T_24_addr = 5'h15;
  assign entries_pte_W__T_24_mask = 1'h0;
  assign entries_pte_W__T_24_en = reset | _T_1;
  assign entries_pte_W__T_25_data = 1'h0;
  assign entries_pte_W__T_25_addr = 5'h16;
  assign entries_pte_W__T_25_mask = 1'h0;
  assign entries_pte_W__T_25_en = reset | _T_1;
  assign entries_pte_W__T_26_data = 1'h0;
  assign entries_pte_W__T_26_addr = 5'h17;
  assign entries_pte_W__T_26_mask = 1'h0;
  assign entries_pte_W__T_26_en = reset | _T_1;
  assign entries_pte_W__T_27_data = 1'h0;
  assign entries_pte_W__T_27_addr = 5'h18;
  assign entries_pte_W__T_27_mask = 1'h0;
  assign entries_pte_W__T_27_en = reset | _T_1;
  assign entries_pte_W__T_28_data = 1'h0;
  assign entries_pte_W__T_28_addr = 5'h19;
  assign entries_pte_W__T_28_mask = 1'h0;
  assign entries_pte_W__T_28_en = reset | _T_1;
  assign entries_pte_W__T_29_data = 1'h0;
  assign entries_pte_W__T_29_addr = 5'h1a;
  assign entries_pte_W__T_29_mask = 1'h0;
  assign entries_pte_W__T_29_en = reset | _T_1;
  assign entries_pte_W__T_30_data = 1'h0;
  assign entries_pte_W__T_30_addr = 5'h1b;
  assign entries_pte_W__T_30_mask = 1'h0;
  assign entries_pte_W__T_30_en = reset | _T_1;
  assign entries_pte_W__T_31_data = 1'h0;
  assign entries_pte_W__T_31_addr = 5'h1c;
  assign entries_pte_W__T_31_mask = 1'h0;
  assign entries_pte_W__T_31_en = reset | _T_1;
  assign entries_pte_W__T_32_data = 1'h0;
  assign entries_pte_W__T_32_addr = 5'h1d;
  assign entries_pte_W__T_32_mask = 1'h0;
  assign entries_pte_W__T_32_en = reset | _T_1;
  assign entries_pte_W__T_33_data = 1'h0;
  assign entries_pte_W__T_33_addr = 5'h1e;
  assign entries_pte_W__T_33_mask = 1'h0;
  assign entries_pte_W__T_33_en = reset | _T_1;
  assign entries_pte_W__T_34_data = 1'h0;
  assign entries_pte_W__T_34_addr = 5'h1f;
  assign entries_pte_W__T_34_mask = 1'h0;
  assign entries_pte_W__T_34_en = reset | _T_1;
  assign entries_pte_W__T_57_data = 1'h0;
  assign entries_pte_W__T_57_addr = _T_55[4:0];
  assign entries_pte_W__T_57_mask = 1'h0;
  assign entries_pte_W__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_W__T_58_data = 1'h0;
  assign entries_pte_W__T_58_addr = _T_55[4:0];
  assign entries_pte_W__T_58_mask = 1'h0;
  assign entries_pte_W__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_W__T_59_data = io_modify_pte_W;
  assign entries_pte_W__T_59_addr = _T_55[4:0];
  assign entries_pte_W__T_59_mask = 1'h1;
  assign entries_pte_W__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_W__T_65_data = 1'h0;
  assign entries_pte_W__T_65_addr = _T_55[4:0];
  assign entries_pte_W__T_65_mask = 1'h0;
  assign entries_pte_W__T_65_en = _T_60 & _T_64;
  assign entries_pte_R__T_39_addr = _T_37[4:0];
  assign entries_pte_R__T_39_data = entries_pte_R[entries_pte_R__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_R__T_49_addr = _T_47[4:0];
  assign entries_pte_R__T_49_data = entries_pte_R[entries_pte_R__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_R__T_61_addr = _T_55[4:0];
  assign entries_pte_R__T_61_data = entries_pte_R[entries_pte_R__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_R__T_3_data = 1'h0;
  assign entries_pte_R__T_3_addr = 5'h0;
  assign entries_pte_R__T_3_mask = 1'h0;
  assign entries_pte_R__T_3_en = reset | _T_1;
  assign entries_pte_R__T_4_data = 1'h0;
  assign entries_pte_R__T_4_addr = 5'h1;
  assign entries_pte_R__T_4_mask = 1'h0;
  assign entries_pte_R__T_4_en = reset | _T_1;
  assign entries_pte_R__T_5_data = 1'h0;
  assign entries_pte_R__T_5_addr = 5'h2;
  assign entries_pte_R__T_5_mask = 1'h0;
  assign entries_pte_R__T_5_en = reset | _T_1;
  assign entries_pte_R__T_6_data = 1'h0;
  assign entries_pte_R__T_6_addr = 5'h3;
  assign entries_pte_R__T_6_mask = 1'h0;
  assign entries_pte_R__T_6_en = reset | _T_1;
  assign entries_pte_R__T_7_data = 1'h0;
  assign entries_pte_R__T_7_addr = 5'h4;
  assign entries_pte_R__T_7_mask = 1'h0;
  assign entries_pte_R__T_7_en = reset | _T_1;
  assign entries_pte_R__T_8_data = 1'h0;
  assign entries_pte_R__T_8_addr = 5'h5;
  assign entries_pte_R__T_8_mask = 1'h0;
  assign entries_pte_R__T_8_en = reset | _T_1;
  assign entries_pte_R__T_9_data = 1'h0;
  assign entries_pte_R__T_9_addr = 5'h6;
  assign entries_pte_R__T_9_mask = 1'h0;
  assign entries_pte_R__T_9_en = reset | _T_1;
  assign entries_pte_R__T_10_data = 1'h0;
  assign entries_pte_R__T_10_addr = 5'h7;
  assign entries_pte_R__T_10_mask = 1'h0;
  assign entries_pte_R__T_10_en = reset | _T_1;
  assign entries_pte_R__T_11_data = 1'h0;
  assign entries_pte_R__T_11_addr = 5'h8;
  assign entries_pte_R__T_11_mask = 1'h0;
  assign entries_pte_R__T_11_en = reset | _T_1;
  assign entries_pte_R__T_12_data = 1'h0;
  assign entries_pte_R__T_12_addr = 5'h9;
  assign entries_pte_R__T_12_mask = 1'h0;
  assign entries_pte_R__T_12_en = reset | _T_1;
  assign entries_pte_R__T_13_data = 1'h0;
  assign entries_pte_R__T_13_addr = 5'ha;
  assign entries_pte_R__T_13_mask = 1'h0;
  assign entries_pte_R__T_13_en = reset | _T_1;
  assign entries_pte_R__T_14_data = 1'h0;
  assign entries_pte_R__T_14_addr = 5'hb;
  assign entries_pte_R__T_14_mask = 1'h0;
  assign entries_pte_R__T_14_en = reset | _T_1;
  assign entries_pte_R__T_15_data = 1'h0;
  assign entries_pte_R__T_15_addr = 5'hc;
  assign entries_pte_R__T_15_mask = 1'h0;
  assign entries_pte_R__T_15_en = reset | _T_1;
  assign entries_pte_R__T_16_data = 1'h0;
  assign entries_pte_R__T_16_addr = 5'hd;
  assign entries_pte_R__T_16_mask = 1'h0;
  assign entries_pte_R__T_16_en = reset | _T_1;
  assign entries_pte_R__T_17_data = 1'h0;
  assign entries_pte_R__T_17_addr = 5'he;
  assign entries_pte_R__T_17_mask = 1'h0;
  assign entries_pte_R__T_17_en = reset | _T_1;
  assign entries_pte_R__T_18_data = 1'h0;
  assign entries_pte_R__T_18_addr = 5'hf;
  assign entries_pte_R__T_18_mask = 1'h0;
  assign entries_pte_R__T_18_en = reset | _T_1;
  assign entries_pte_R__T_19_data = 1'h0;
  assign entries_pte_R__T_19_addr = 5'h10;
  assign entries_pte_R__T_19_mask = 1'h0;
  assign entries_pte_R__T_19_en = reset | _T_1;
  assign entries_pte_R__T_20_data = 1'h0;
  assign entries_pte_R__T_20_addr = 5'h11;
  assign entries_pte_R__T_20_mask = 1'h0;
  assign entries_pte_R__T_20_en = reset | _T_1;
  assign entries_pte_R__T_21_data = 1'h0;
  assign entries_pte_R__T_21_addr = 5'h12;
  assign entries_pte_R__T_21_mask = 1'h0;
  assign entries_pte_R__T_21_en = reset | _T_1;
  assign entries_pte_R__T_22_data = 1'h0;
  assign entries_pte_R__T_22_addr = 5'h13;
  assign entries_pte_R__T_22_mask = 1'h0;
  assign entries_pte_R__T_22_en = reset | _T_1;
  assign entries_pte_R__T_23_data = 1'h0;
  assign entries_pte_R__T_23_addr = 5'h14;
  assign entries_pte_R__T_23_mask = 1'h0;
  assign entries_pte_R__T_23_en = reset | _T_1;
  assign entries_pte_R__T_24_data = 1'h0;
  assign entries_pte_R__T_24_addr = 5'h15;
  assign entries_pte_R__T_24_mask = 1'h0;
  assign entries_pte_R__T_24_en = reset | _T_1;
  assign entries_pte_R__T_25_data = 1'h0;
  assign entries_pte_R__T_25_addr = 5'h16;
  assign entries_pte_R__T_25_mask = 1'h0;
  assign entries_pte_R__T_25_en = reset | _T_1;
  assign entries_pte_R__T_26_data = 1'h0;
  assign entries_pte_R__T_26_addr = 5'h17;
  assign entries_pte_R__T_26_mask = 1'h0;
  assign entries_pte_R__T_26_en = reset | _T_1;
  assign entries_pte_R__T_27_data = 1'h0;
  assign entries_pte_R__T_27_addr = 5'h18;
  assign entries_pte_R__T_27_mask = 1'h0;
  assign entries_pte_R__T_27_en = reset | _T_1;
  assign entries_pte_R__T_28_data = 1'h0;
  assign entries_pte_R__T_28_addr = 5'h19;
  assign entries_pte_R__T_28_mask = 1'h0;
  assign entries_pte_R__T_28_en = reset | _T_1;
  assign entries_pte_R__T_29_data = 1'h0;
  assign entries_pte_R__T_29_addr = 5'h1a;
  assign entries_pte_R__T_29_mask = 1'h0;
  assign entries_pte_R__T_29_en = reset | _T_1;
  assign entries_pte_R__T_30_data = 1'h0;
  assign entries_pte_R__T_30_addr = 5'h1b;
  assign entries_pte_R__T_30_mask = 1'h0;
  assign entries_pte_R__T_30_en = reset | _T_1;
  assign entries_pte_R__T_31_data = 1'h0;
  assign entries_pte_R__T_31_addr = 5'h1c;
  assign entries_pte_R__T_31_mask = 1'h0;
  assign entries_pte_R__T_31_en = reset | _T_1;
  assign entries_pte_R__T_32_data = 1'h0;
  assign entries_pte_R__T_32_addr = 5'h1d;
  assign entries_pte_R__T_32_mask = 1'h0;
  assign entries_pte_R__T_32_en = reset | _T_1;
  assign entries_pte_R__T_33_data = 1'h0;
  assign entries_pte_R__T_33_addr = 5'h1e;
  assign entries_pte_R__T_33_mask = 1'h0;
  assign entries_pte_R__T_33_en = reset | _T_1;
  assign entries_pte_R__T_34_data = 1'h0;
  assign entries_pte_R__T_34_addr = 5'h1f;
  assign entries_pte_R__T_34_mask = 1'h0;
  assign entries_pte_R__T_34_en = reset | _T_1;
  assign entries_pte_R__T_57_data = 1'h0;
  assign entries_pte_R__T_57_addr = _T_55[4:0];
  assign entries_pte_R__T_57_mask = 1'h0;
  assign entries_pte_R__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_R__T_58_data = 1'h0;
  assign entries_pte_R__T_58_addr = _T_55[4:0];
  assign entries_pte_R__T_58_mask = 1'h0;
  assign entries_pte_R__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_R__T_59_data = io_modify_pte_R;
  assign entries_pte_R__T_59_addr = _T_55[4:0];
  assign entries_pte_R__T_59_mask = 1'h1;
  assign entries_pte_R__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_R__T_65_data = 1'h0;
  assign entries_pte_R__T_65_addr = _T_55[4:0];
  assign entries_pte_R__T_65_mask = 1'h0;
  assign entries_pte_R__T_65_en = _T_60 & _T_64;
  assign entries_pte_V__T_39_addr = _T_37[4:0];
  assign entries_pte_V__T_39_data = entries_pte_V[entries_pte_V__T_39_addr]; // @[TLB.scala 38:20]
  assign entries_pte_V__T_49_addr = _T_47[4:0];
  assign entries_pte_V__T_49_data = entries_pte_V[entries_pte_V__T_49_addr]; // @[TLB.scala 38:20]
  assign entries_pte_V__T_61_addr = _T_55[4:0];
  assign entries_pte_V__T_61_data = entries_pte_V[entries_pte_V__T_61_addr]; // @[TLB.scala 38:20]
  assign entries_pte_V__T_3_data = 1'h0;
  assign entries_pte_V__T_3_addr = 5'h0;
  assign entries_pte_V__T_3_mask = 1'h0;
  assign entries_pte_V__T_3_en = reset | _T_1;
  assign entries_pte_V__T_4_data = 1'h0;
  assign entries_pte_V__T_4_addr = 5'h1;
  assign entries_pte_V__T_4_mask = 1'h0;
  assign entries_pte_V__T_4_en = reset | _T_1;
  assign entries_pte_V__T_5_data = 1'h0;
  assign entries_pte_V__T_5_addr = 5'h2;
  assign entries_pte_V__T_5_mask = 1'h0;
  assign entries_pte_V__T_5_en = reset | _T_1;
  assign entries_pte_V__T_6_data = 1'h0;
  assign entries_pte_V__T_6_addr = 5'h3;
  assign entries_pte_V__T_6_mask = 1'h0;
  assign entries_pte_V__T_6_en = reset | _T_1;
  assign entries_pte_V__T_7_data = 1'h0;
  assign entries_pte_V__T_7_addr = 5'h4;
  assign entries_pte_V__T_7_mask = 1'h0;
  assign entries_pte_V__T_7_en = reset | _T_1;
  assign entries_pte_V__T_8_data = 1'h0;
  assign entries_pte_V__T_8_addr = 5'h5;
  assign entries_pte_V__T_8_mask = 1'h0;
  assign entries_pte_V__T_8_en = reset | _T_1;
  assign entries_pte_V__T_9_data = 1'h0;
  assign entries_pte_V__T_9_addr = 5'h6;
  assign entries_pte_V__T_9_mask = 1'h0;
  assign entries_pte_V__T_9_en = reset | _T_1;
  assign entries_pte_V__T_10_data = 1'h0;
  assign entries_pte_V__T_10_addr = 5'h7;
  assign entries_pte_V__T_10_mask = 1'h0;
  assign entries_pte_V__T_10_en = reset | _T_1;
  assign entries_pte_V__T_11_data = 1'h0;
  assign entries_pte_V__T_11_addr = 5'h8;
  assign entries_pte_V__T_11_mask = 1'h0;
  assign entries_pte_V__T_11_en = reset | _T_1;
  assign entries_pte_V__T_12_data = 1'h0;
  assign entries_pte_V__T_12_addr = 5'h9;
  assign entries_pte_V__T_12_mask = 1'h0;
  assign entries_pte_V__T_12_en = reset | _T_1;
  assign entries_pte_V__T_13_data = 1'h0;
  assign entries_pte_V__T_13_addr = 5'ha;
  assign entries_pte_V__T_13_mask = 1'h0;
  assign entries_pte_V__T_13_en = reset | _T_1;
  assign entries_pte_V__T_14_data = 1'h0;
  assign entries_pte_V__T_14_addr = 5'hb;
  assign entries_pte_V__T_14_mask = 1'h0;
  assign entries_pte_V__T_14_en = reset | _T_1;
  assign entries_pte_V__T_15_data = 1'h0;
  assign entries_pte_V__T_15_addr = 5'hc;
  assign entries_pte_V__T_15_mask = 1'h0;
  assign entries_pte_V__T_15_en = reset | _T_1;
  assign entries_pte_V__T_16_data = 1'h0;
  assign entries_pte_V__T_16_addr = 5'hd;
  assign entries_pte_V__T_16_mask = 1'h0;
  assign entries_pte_V__T_16_en = reset | _T_1;
  assign entries_pte_V__T_17_data = 1'h0;
  assign entries_pte_V__T_17_addr = 5'he;
  assign entries_pte_V__T_17_mask = 1'h0;
  assign entries_pte_V__T_17_en = reset | _T_1;
  assign entries_pte_V__T_18_data = 1'h0;
  assign entries_pte_V__T_18_addr = 5'hf;
  assign entries_pte_V__T_18_mask = 1'h0;
  assign entries_pte_V__T_18_en = reset | _T_1;
  assign entries_pte_V__T_19_data = 1'h0;
  assign entries_pte_V__T_19_addr = 5'h10;
  assign entries_pte_V__T_19_mask = 1'h0;
  assign entries_pte_V__T_19_en = reset | _T_1;
  assign entries_pte_V__T_20_data = 1'h0;
  assign entries_pte_V__T_20_addr = 5'h11;
  assign entries_pte_V__T_20_mask = 1'h0;
  assign entries_pte_V__T_20_en = reset | _T_1;
  assign entries_pte_V__T_21_data = 1'h0;
  assign entries_pte_V__T_21_addr = 5'h12;
  assign entries_pte_V__T_21_mask = 1'h0;
  assign entries_pte_V__T_21_en = reset | _T_1;
  assign entries_pte_V__T_22_data = 1'h0;
  assign entries_pte_V__T_22_addr = 5'h13;
  assign entries_pte_V__T_22_mask = 1'h0;
  assign entries_pte_V__T_22_en = reset | _T_1;
  assign entries_pte_V__T_23_data = 1'h0;
  assign entries_pte_V__T_23_addr = 5'h14;
  assign entries_pte_V__T_23_mask = 1'h0;
  assign entries_pte_V__T_23_en = reset | _T_1;
  assign entries_pte_V__T_24_data = 1'h0;
  assign entries_pte_V__T_24_addr = 5'h15;
  assign entries_pte_V__T_24_mask = 1'h0;
  assign entries_pte_V__T_24_en = reset | _T_1;
  assign entries_pte_V__T_25_data = 1'h0;
  assign entries_pte_V__T_25_addr = 5'h16;
  assign entries_pte_V__T_25_mask = 1'h0;
  assign entries_pte_V__T_25_en = reset | _T_1;
  assign entries_pte_V__T_26_data = 1'h0;
  assign entries_pte_V__T_26_addr = 5'h17;
  assign entries_pte_V__T_26_mask = 1'h0;
  assign entries_pte_V__T_26_en = reset | _T_1;
  assign entries_pte_V__T_27_data = 1'h0;
  assign entries_pte_V__T_27_addr = 5'h18;
  assign entries_pte_V__T_27_mask = 1'h0;
  assign entries_pte_V__T_27_en = reset | _T_1;
  assign entries_pte_V__T_28_data = 1'h0;
  assign entries_pte_V__T_28_addr = 5'h19;
  assign entries_pte_V__T_28_mask = 1'h0;
  assign entries_pte_V__T_28_en = reset | _T_1;
  assign entries_pte_V__T_29_data = 1'h0;
  assign entries_pte_V__T_29_addr = 5'h1a;
  assign entries_pte_V__T_29_mask = 1'h0;
  assign entries_pte_V__T_29_en = reset | _T_1;
  assign entries_pte_V__T_30_data = 1'h0;
  assign entries_pte_V__T_30_addr = 5'h1b;
  assign entries_pte_V__T_30_mask = 1'h0;
  assign entries_pte_V__T_30_en = reset | _T_1;
  assign entries_pte_V__T_31_data = 1'h0;
  assign entries_pte_V__T_31_addr = 5'h1c;
  assign entries_pte_V__T_31_mask = 1'h0;
  assign entries_pte_V__T_31_en = reset | _T_1;
  assign entries_pte_V__T_32_data = 1'h0;
  assign entries_pte_V__T_32_addr = 5'h1d;
  assign entries_pte_V__T_32_mask = 1'h0;
  assign entries_pte_V__T_32_en = reset | _T_1;
  assign entries_pte_V__T_33_data = 1'h0;
  assign entries_pte_V__T_33_addr = 5'h1e;
  assign entries_pte_V__T_33_mask = 1'h0;
  assign entries_pte_V__T_33_en = reset | _T_1;
  assign entries_pte_V__T_34_data = 1'h0;
  assign entries_pte_V__T_34_addr = 5'h1f;
  assign entries_pte_V__T_34_mask = 1'h0;
  assign entries_pte_V__T_34_en = reset | _T_1;
  assign entries_pte_V__T_57_data = 1'h0;
  assign entries_pte_V__T_57_addr = _T_55[4:0];
  assign entries_pte_V__T_57_mask = 1'h0;
  assign entries_pte_V__T_57_en = io_modify_mode == 2'h1;
  assign entries_pte_V__T_58_data = 1'h0;
  assign entries_pte_V__T_58_addr = _T_55[4:0];
  assign entries_pte_V__T_58_mask = 1'h0;
  assign entries_pte_V__T_58_en = io_modify_mode == 2'h1;
  assign entries_pte_V__T_59_data = io_modify_pte_V;
  assign entries_pte_V__T_59_addr = _T_55[4:0];
  assign entries_pte_V__T_59_mask = 1'h1;
  assign entries_pte_V__T_59_en = io_modify_mode == 2'h1;
  assign entries_pte_V__T_65_data = 1'h0;
  assign entries_pte_V__T_65_addr = _T_55[4:0];
  assign entries_pte_V__T_65_mask = 1'h0;
  assign entries_pte_V__T_65_en = _T_60 & _T_64;
  assign io_query_rsp_valid = reset ? io_query_req_valid : _T_44; // @[TLB.scala 56:19 TLB.scala 67:19]
  assign io_query_rsp_bits_ppn_p2 = reset ? io_query_req_bits_p2 : entries_pte_ppn_p2__T_39_data; // @[TLB.scala 57:18 TLB.scala 58:22 TLB.scala 68:18]
  assign io_query_rsp_bits_ppn_p1 = reset ? io_query_req_bits_p1 : entries_pte_ppn_p1__T_39_data; // @[TLB.scala 57:18 TLB.scala 58:22 TLB.scala 68:18]
  assign io_query_rsp_bits_U = reset | entries_pte_U__T_39_data; // @[TLB.scala 57:18 TLB.scala 63:20 TLB.scala 68:18]
  assign io_query_rsp_bits_X = reset | entries_pte_X__T_39_data; // @[TLB.scala 57:18 TLB.scala 60:20 TLB.scala 68:18]
  assign io_query_rsp_bits_V = reset | entries_pte_V__T_39_data; // @[TLB.scala 57:18 TLB.scala 59:20 TLB.scala 68:18]
  assign io_query2_rsp_valid = reset ? io_query2_req_valid : _T_54; // @[TLB.scala 56:19 TLB.scala 67:19]
  assign io_query2_rsp_bits_ppn_p2 = reset ? io_query2_req_bits_p2 : entries_pte_ppn_p2__T_49_data; // @[TLB.scala 57:18 TLB.scala 58:22 TLB.scala 68:18]
  assign io_query2_rsp_bits_ppn_p1 = reset ? io_query2_req_bits_p1 : entries_pte_ppn_p1__T_49_data; // @[TLB.scala 57:18 TLB.scala 58:22 TLB.scala 68:18]
  assign io_query2_rsp_bits_U = reset | entries_pte_U__T_49_data; // @[TLB.scala 57:18 TLB.scala 63:20 TLB.scala 68:18]
  assign io_query2_rsp_bits_X = reset | entries_pte_X__T_49_data; // @[TLB.scala 57:18 TLB.scala 60:20 TLB.scala 68:18]
  assign io_query2_rsp_bits_W = reset | entries_pte_W__T_49_data; // @[TLB.scala 57:18 TLB.scala 62:20 TLB.scala 68:18]
  assign io_query2_rsp_bits_R = reset | entries_pte_R__T_49_data; // @[TLB.scala 57:18 TLB.scala 61:20 TLB.scala 68:18]
  assign io_query2_rsp_bits_V = reset | entries_pte_V__T_49_data; // @[TLB.scala 57:18 TLB.scala 59:20 TLB.scala 68:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_valid[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_vpn_p2[initvar] = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_vpn_p1[initvar] = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_ppn_p2[initvar] = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_ppn_p1[initvar] = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_U[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_X[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_W[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_R[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    entries_pte_V[initvar] = _RAND_9[0:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(entries_valid__T_3_en & entries_valid__T_3_mask) begin
      entries_valid[entries_valid__T_3_addr] <= entries_valid__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_4_en & entries_valid__T_4_mask) begin
      entries_valid[entries_valid__T_4_addr] <= entries_valid__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_5_en & entries_valid__T_5_mask) begin
      entries_valid[entries_valid__T_5_addr] <= entries_valid__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_6_en & entries_valid__T_6_mask) begin
      entries_valid[entries_valid__T_6_addr] <= entries_valid__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_7_en & entries_valid__T_7_mask) begin
      entries_valid[entries_valid__T_7_addr] <= entries_valid__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_8_en & entries_valid__T_8_mask) begin
      entries_valid[entries_valid__T_8_addr] <= entries_valid__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_9_en & entries_valid__T_9_mask) begin
      entries_valid[entries_valid__T_9_addr] <= entries_valid__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_10_en & entries_valid__T_10_mask) begin
      entries_valid[entries_valid__T_10_addr] <= entries_valid__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_11_en & entries_valid__T_11_mask) begin
      entries_valid[entries_valid__T_11_addr] <= entries_valid__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_12_en & entries_valid__T_12_mask) begin
      entries_valid[entries_valid__T_12_addr] <= entries_valid__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_13_en & entries_valid__T_13_mask) begin
      entries_valid[entries_valid__T_13_addr] <= entries_valid__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_14_en & entries_valid__T_14_mask) begin
      entries_valid[entries_valid__T_14_addr] <= entries_valid__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_15_en & entries_valid__T_15_mask) begin
      entries_valid[entries_valid__T_15_addr] <= entries_valid__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_16_en & entries_valid__T_16_mask) begin
      entries_valid[entries_valid__T_16_addr] <= entries_valid__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_17_en & entries_valid__T_17_mask) begin
      entries_valid[entries_valid__T_17_addr] <= entries_valid__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_18_en & entries_valid__T_18_mask) begin
      entries_valid[entries_valid__T_18_addr] <= entries_valid__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_19_en & entries_valid__T_19_mask) begin
      entries_valid[entries_valid__T_19_addr] <= entries_valid__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_20_en & entries_valid__T_20_mask) begin
      entries_valid[entries_valid__T_20_addr] <= entries_valid__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_21_en & entries_valid__T_21_mask) begin
      entries_valid[entries_valid__T_21_addr] <= entries_valid__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_22_en & entries_valid__T_22_mask) begin
      entries_valid[entries_valid__T_22_addr] <= entries_valid__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_23_en & entries_valid__T_23_mask) begin
      entries_valid[entries_valid__T_23_addr] <= entries_valid__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_24_en & entries_valid__T_24_mask) begin
      entries_valid[entries_valid__T_24_addr] <= entries_valid__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_25_en & entries_valid__T_25_mask) begin
      entries_valid[entries_valid__T_25_addr] <= entries_valid__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_26_en & entries_valid__T_26_mask) begin
      entries_valid[entries_valid__T_26_addr] <= entries_valid__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_27_en & entries_valid__T_27_mask) begin
      entries_valid[entries_valid__T_27_addr] <= entries_valid__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_28_en & entries_valid__T_28_mask) begin
      entries_valid[entries_valid__T_28_addr] <= entries_valid__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_29_en & entries_valid__T_29_mask) begin
      entries_valid[entries_valid__T_29_addr] <= entries_valid__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_30_en & entries_valid__T_30_mask) begin
      entries_valid[entries_valid__T_30_addr] <= entries_valid__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_31_en & entries_valid__T_31_mask) begin
      entries_valid[entries_valid__T_31_addr] <= entries_valid__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_32_en & entries_valid__T_32_mask) begin
      entries_valid[entries_valid__T_32_addr] <= entries_valid__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_33_en & entries_valid__T_33_mask) begin
      entries_valid[entries_valid__T_33_addr] <= entries_valid__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_34_en & entries_valid__T_34_mask) begin
      entries_valid[entries_valid__T_34_addr] <= entries_valid__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_57_en & entries_valid__T_57_mask) begin
      entries_valid[entries_valid__T_57_addr] <= entries_valid__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_58_en & entries_valid__T_58_mask) begin
      entries_valid[entries_valid__T_58_addr] <= entries_valid__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_59_en & entries_valid__T_59_mask) begin
      entries_valid[entries_valid__T_59_addr] <= entries_valid__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_valid__T_65_en & entries_valid__T_65_mask) begin
      entries_valid[entries_valid__T_65_addr] <= entries_valid__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_3_en & entries_vpn_p2__T_3_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_3_addr] <= entries_vpn_p2__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_4_en & entries_vpn_p2__T_4_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_4_addr] <= entries_vpn_p2__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_5_en & entries_vpn_p2__T_5_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_5_addr] <= entries_vpn_p2__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_6_en & entries_vpn_p2__T_6_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_6_addr] <= entries_vpn_p2__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_7_en & entries_vpn_p2__T_7_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_7_addr] <= entries_vpn_p2__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_8_en & entries_vpn_p2__T_8_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_8_addr] <= entries_vpn_p2__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_9_en & entries_vpn_p2__T_9_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_9_addr] <= entries_vpn_p2__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_10_en & entries_vpn_p2__T_10_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_10_addr] <= entries_vpn_p2__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_11_en & entries_vpn_p2__T_11_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_11_addr] <= entries_vpn_p2__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_12_en & entries_vpn_p2__T_12_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_12_addr] <= entries_vpn_p2__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_13_en & entries_vpn_p2__T_13_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_13_addr] <= entries_vpn_p2__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_14_en & entries_vpn_p2__T_14_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_14_addr] <= entries_vpn_p2__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_15_en & entries_vpn_p2__T_15_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_15_addr] <= entries_vpn_p2__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_16_en & entries_vpn_p2__T_16_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_16_addr] <= entries_vpn_p2__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_17_en & entries_vpn_p2__T_17_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_17_addr] <= entries_vpn_p2__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_18_en & entries_vpn_p2__T_18_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_18_addr] <= entries_vpn_p2__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_19_en & entries_vpn_p2__T_19_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_19_addr] <= entries_vpn_p2__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_20_en & entries_vpn_p2__T_20_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_20_addr] <= entries_vpn_p2__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_21_en & entries_vpn_p2__T_21_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_21_addr] <= entries_vpn_p2__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_22_en & entries_vpn_p2__T_22_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_22_addr] <= entries_vpn_p2__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_23_en & entries_vpn_p2__T_23_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_23_addr] <= entries_vpn_p2__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_24_en & entries_vpn_p2__T_24_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_24_addr] <= entries_vpn_p2__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_25_en & entries_vpn_p2__T_25_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_25_addr] <= entries_vpn_p2__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_26_en & entries_vpn_p2__T_26_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_26_addr] <= entries_vpn_p2__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_27_en & entries_vpn_p2__T_27_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_27_addr] <= entries_vpn_p2__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_28_en & entries_vpn_p2__T_28_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_28_addr] <= entries_vpn_p2__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_29_en & entries_vpn_p2__T_29_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_29_addr] <= entries_vpn_p2__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_30_en & entries_vpn_p2__T_30_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_30_addr] <= entries_vpn_p2__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_31_en & entries_vpn_p2__T_31_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_31_addr] <= entries_vpn_p2__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_32_en & entries_vpn_p2__T_32_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_32_addr] <= entries_vpn_p2__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_33_en & entries_vpn_p2__T_33_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_33_addr] <= entries_vpn_p2__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_34_en & entries_vpn_p2__T_34_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_34_addr] <= entries_vpn_p2__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_57_en & entries_vpn_p2__T_57_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_57_addr] <= entries_vpn_p2__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_58_en & entries_vpn_p2__T_58_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_58_addr] <= entries_vpn_p2__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_59_en & entries_vpn_p2__T_59_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_59_addr] <= entries_vpn_p2__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p2__T_65_en & entries_vpn_p2__T_65_mask) begin
      entries_vpn_p2[entries_vpn_p2__T_65_addr] <= entries_vpn_p2__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_3_en & entries_vpn_p1__T_3_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_3_addr] <= entries_vpn_p1__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_4_en & entries_vpn_p1__T_4_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_4_addr] <= entries_vpn_p1__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_5_en & entries_vpn_p1__T_5_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_5_addr] <= entries_vpn_p1__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_6_en & entries_vpn_p1__T_6_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_6_addr] <= entries_vpn_p1__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_7_en & entries_vpn_p1__T_7_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_7_addr] <= entries_vpn_p1__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_8_en & entries_vpn_p1__T_8_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_8_addr] <= entries_vpn_p1__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_9_en & entries_vpn_p1__T_9_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_9_addr] <= entries_vpn_p1__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_10_en & entries_vpn_p1__T_10_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_10_addr] <= entries_vpn_p1__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_11_en & entries_vpn_p1__T_11_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_11_addr] <= entries_vpn_p1__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_12_en & entries_vpn_p1__T_12_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_12_addr] <= entries_vpn_p1__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_13_en & entries_vpn_p1__T_13_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_13_addr] <= entries_vpn_p1__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_14_en & entries_vpn_p1__T_14_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_14_addr] <= entries_vpn_p1__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_15_en & entries_vpn_p1__T_15_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_15_addr] <= entries_vpn_p1__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_16_en & entries_vpn_p1__T_16_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_16_addr] <= entries_vpn_p1__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_17_en & entries_vpn_p1__T_17_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_17_addr] <= entries_vpn_p1__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_18_en & entries_vpn_p1__T_18_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_18_addr] <= entries_vpn_p1__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_19_en & entries_vpn_p1__T_19_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_19_addr] <= entries_vpn_p1__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_20_en & entries_vpn_p1__T_20_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_20_addr] <= entries_vpn_p1__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_21_en & entries_vpn_p1__T_21_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_21_addr] <= entries_vpn_p1__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_22_en & entries_vpn_p1__T_22_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_22_addr] <= entries_vpn_p1__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_23_en & entries_vpn_p1__T_23_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_23_addr] <= entries_vpn_p1__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_24_en & entries_vpn_p1__T_24_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_24_addr] <= entries_vpn_p1__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_25_en & entries_vpn_p1__T_25_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_25_addr] <= entries_vpn_p1__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_26_en & entries_vpn_p1__T_26_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_26_addr] <= entries_vpn_p1__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_27_en & entries_vpn_p1__T_27_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_27_addr] <= entries_vpn_p1__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_28_en & entries_vpn_p1__T_28_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_28_addr] <= entries_vpn_p1__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_29_en & entries_vpn_p1__T_29_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_29_addr] <= entries_vpn_p1__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_30_en & entries_vpn_p1__T_30_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_30_addr] <= entries_vpn_p1__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_31_en & entries_vpn_p1__T_31_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_31_addr] <= entries_vpn_p1__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_32_en & entries_vpn_p1__T_32_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_32_addr] <= entries_vpn_p1__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_33_en & entries_vpn_p1__T_33_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_33_addr] <= entries_vpn_p1__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_34_en & entries_vpn_p1__T_34_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_34_addr] <= entries_vpn_p1__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_57_en & entries_vpn_p1__T_57_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_57_addr] <= entries_vpn_p1__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_58_en & entries_vpn_p1__T_58_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_58_addr] <= entries_vpn_p1__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_59_en & entries_vpn_p1__T_59_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_59_addr] <= entries_vpn_p1__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_vpn_p1__T_65_en & entries_vpn_p1__T_65_mask) begin
      entries_vpn_p1[entries_vpn_p1__T_65_addr] <= entries_vpn_p1__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_3_en & entries_pte_ppn_p2__T_3_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_3_addr] <= entries_pte_ppn_p2__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_4_en & entries_pte_ppn_p2__T_4_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_4_addr] <= entries_pte_ppn_p2__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_5_en & entries_pte_ppn_p2__T_5_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_5_addr] <= entries_pte_ppn_p2__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_6_en & entries_pte_ppn_p2__T_6_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_6_addr] <= entries_pte_ppn_p2__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_7_en & entries_pte_ppn_p2__T_7_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_7_addr] <= entries_pte_ppn_p2__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_8_en & entries_pte_ppn_p2__T_8_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_8_addr] <= entries_pte_ppn_p2__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_9_en & entries_pte_ppn_p2__T_9_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_9_addr] <= entries_pte_ppn_p2__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_10_en & entries_pte_ppn_p2__T_10_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_10_addr] <= entries_pte_ppn_p2__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_11_en & entries_pte_ppn_p2__T_11_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_11_addr] <= entries_pte_ppn_p2__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_12_en & entries_pte_ppn_p2__T_12_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_12_addr] <= entries_pte_ppn_p2__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_13_en & entries_pte_ppn_p2__T_13_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_13_addr] <= entries_pte_ppn_p2__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_14_en & entries_pte_ppn_p2__T_14_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_14_addr] <= entries_pte_ppn_p2__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_15_en & entries_pte_ppn_p2__T_15_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_15_addr] <= entries_pte_ppn_p2__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_16_en & entries_pte_ppn_p2__T_16_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_16_addr] <= entries_pte_ppn_p2__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_17_en & entries_pte_ppn_p2__T_17_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_17_addr] <= entries_pte_ppn_p2__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_18_en & entries_pte_ppn_p2__T_18_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_18_addr] <= entries_pte_ppn_p2__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_19_en & entries_pte_ppn_p2__T_19_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_19_addr] <= entries_pte_ppn_p2__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_20_en & entries_pte_ppn_p2__T_20_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_20_addr] <= entries_pte_ppn_p2__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_21_en & entries_pte_ppn_p2__T_21_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_21_addr] <= entries_pte_ppn_p2__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_22_en & entries_pte_ppn_p2__T_22_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_22_addr] <= entries_pte_ppn_p2__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_23_en & entries_pte_ppn_p2__T_23_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_23_addr] <= entries_pte_ppn_p2__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_24_en & entries_pte_ppn_p2__T_24_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_24_addr] <= entries_pte_ppn_p2__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_25_en & entries_pte_ppn_p2__T_25_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_25_addr] <= entries_pte_ppn_p2__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_26_en & entries_pte_ppn_p2__T_26_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_26_addr] <= entries_pte_ppn_p2__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_27_en & entries_pte_ppn_p2__T_27_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_27_addr] <= entries_pte_ppn_p2__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_28_en & entries_pte_ppn_p2__T_28_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_28_addr] <= entries_pte_ppn_p2__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_29_en & entries_pte_ppn_p2__T_29_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_29_addr] <= entries_pte_ppn_p2__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_30_en & entries_pte_ppn_p2__T_30_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_30_addr] <= entries_pte_ppn_p2__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_31_en & entries_pte_ppn_p2__T_31_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_31_addr] <= entries_pte_ppn_p2__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_32_en & entries_pte_ppn_p2__T_32_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_32_addr] <= entries_pte_ppn_p2__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_33_en & entries_pte_ppn_p2__T_33_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_33_addr] <= entries_pte_ppn_p2__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_34_en & entries_pte_ppn_p2__T_34_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_34_addr] <= entries_pte_ppn_p2__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_57_en & entries_pte_ppn_p2__T_57_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_57_addr] <= entries_pte_ppn_p2__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_58_en & entries_pte_ppn_p2__T_58_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_58_addr] <= entries_pte_ppn_p2__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_59_en & entries_pte_ppn_p2__T_59_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_59_addr] <= entries_pte_ppn_p2__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p2__T_65_en & entries_pte_ppn_p2__T_65_mask) begin
      entries_pte_ppn_p2[entries_pte_ppn_p2__T_65_addr] <= entries_pte_ppn_p2__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_3_en & entries_pte_ppn_p1__T_3_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_3_addr] <= entries_pte_ppn_p1__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_4_en & entries_pte_ppn_p1__T_4_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_4_addr] <= entries_pte_ppn_p1__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_5_en & entries_pte_ppn_p1__T_5_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_5_addr] <= entries_pte_ppn_p1__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_6_en & entries_pte_ppn_p1__T_6_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_6_addr] <= entries_pte_ppn_p1__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_7_en & entries_pte_ppn_p1__T_7_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_7_addr] <= entries_pte_ppn_p1__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_8_en & entries_pte_ppn_p1__T_8_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_8_addr] <= entries_pte_ppn_p1__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_9_en & entries_pte_ppn_p1__T_9_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_9_addr] <= entries_pte_ppn_p1__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_10_en & entries_pte_ppn_p1__T_10_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_10_addr] <= entries_pte_ppn_p1__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_11_en & entries_pte_ppn_p1__T_11_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_11_addr] <= entries_pte_ppn_p1__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_12_en & entries_pte_ppn_p1__T_12_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_12_addr] <= entries_pte_ppn_p1__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_13_en & entries_pte_ppn_p1__T_13_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_13_addr] <= entries_pte_ppn_p1__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_14_en & entries_pte_ppn_p1__T_14_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_14_addr] <= entries_pte_ppn_p1__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_15_en & entries_pte_ppn_p1__T_15_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_15_addr] <= entries_pte_ppn_p1__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_16_en & entries_pte_ppn_p1__T_16_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_16_addr] <= entries_pte_ppn_p1__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_17_en & entries_pte_ppn_p1__T_17_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_17_addr] <= entries_pte_ppn_p1__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_18_en & entries_pte_ppn_p1__T_18_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_18_addr] <= entries_pte_ppn_p1__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_19_en & entries_pte_ppn_p1__T_19_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_19_addr] <= entries_pte_ppn_p1__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_20_en & entries_pte_ppn_p1__T_20_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_20_addr] <= entries_pte_ppn_p1__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_21_en & entries_pte_ppn_p1__T_21_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_21_addr] <= entries_pte_ppn_p1__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_22_en & entries_pte_ppn_p1__T_22_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_22_addr] <= entries_pte_ppn_p1__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_23_en & entries_pte_ppn_p1__T_23_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_23_addr] <= entries_pte_ppn_p1__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_24_en & entries_pte_ppn_p1__T_24_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_24_addr] <= entries_pte_ppn_p1__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_25_en & entries_pte_ppn_p1__T_25_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_25_addr] <= entries_pte_ppn_p1__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_26_en & entries_pte_ppn_p1__T_26_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_26_addr] <= entries_pte_ppn_p1__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_27_en & entries_pte_ppn_p1__T_27_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_27_addr] <= entries_pte_ppn_p1__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_28_en & entries_pte_ppn_p1__T_28_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_28_addr] <= entries_pte_ppn_p1__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_29_en & entries_pte_ppn_p1__T_29_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_29_addr] <= entries_pte_ppn_p1__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_30_en & entries_pte_ppn_p1__T_30_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_30_addr] <= entries_pte_ppn_p1__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_31_en & entries_pte_ppn_p1__T_31_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_31_addr] <= entries_pte_ppn_p1__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_32_en & entries_pte_ppn_p1__T_32_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_32_addr] <= entries_pte_ppn_p1__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_33_en & entries_pte_ppn_p1__T_33_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_33_addr] <= entries_pte_ppn_p1__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_34_en & entries_pte_ppn_p1__T_34_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_34_addr] <= entries_pte_ppn_p1__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_57_en & entries_pte_ppn_p1__T_57_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_57_addr] <= entries_pte_ppn_p1__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_58_en & entries_pte_ppn_p1__T_58_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_58_addr] <= entries_pte_ppn_p1__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_59_en & entries_pte_ppn_p1__T_59_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_59_addr] <= entries_pte_ppn_p1__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_ppn_p1__T_65_en & entries_pte_ppn_p1__T_65_mask) begin
      entries_pte_ppn_p1[entries_pte_ppn_p1__T_65_addr] <= entries_pte_ppn_p1__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_3_en & entries_pte_U__T_3_mask) begin
      entries_pte_U[entries_pte_U__T_3_addr] <= entries_pte_U__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_4_en & entries_pte_U__T_4_mask) begin
      entries_pte_U[entries_pte_U__T_4_addr] <= entries_pte_U__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_5_en & entries_pte_U__T_5_mask) begin
      entries_pte_U[entries_pte_U__T_5_addr] <= entries_pte_U__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_6_en & entries_pte_U__T_6_mask) begin
      entries_pte_U[entries_pte_U__T_6_addr] <= entries_pte_U__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_7_en & entries_pte_U__T_7_mask) begin
      entries_pte_U[entries_pte_U__T_7_addr] <= entries_pte_U__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_8_en & entries_pte_U__T_8_mask) begin
      entries_pte_U[entries_pte_U__T_8_addr] <= entries_pte_U__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_9_en & entries_pte_U__T_9_mask) begin
      entries_pte_U[entries_pte_U__T_9_addr] <= entries_pte_U__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_10_en & entries_pte_U__T_10_mask) begin
      entries_pte_U[entries_pte_U__T_10_addr] <= entries_pte_U__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_11_en & entries_pte_U__T_11_mask) begin
      entries_pte_U[entries_pte_U__T_11_addr] <= entries_pte_U__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_12_en & entries_pte_U__T_12_mask) begin
      entries_pte_U[entries_pte_U__T_12_addr] <= entries_pte_U__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_13_en & entries_pte_U__T_13_mask) begin
      entries_pte_U[entries_pte_U__T_13_addr] <= entries_pte_U__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_14_en & entries_pte_U__T_14_mask) begin
      entries_pte_U[entries_pte_U__T_14_addr] <= entries_pte_U__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_15_en & entries_pte_U__T_15_mask) begin
      entries_pte_U[entries_pte_U__T_15_addr] <= entries_pte_U__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_16_en & entries_pte_U__T_16_mask) begin
      entries_pte_U[entries_pte_U__T_16_addr] <= entries_pte_U__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_17_en & entries_pte_U__T_17_mask) begin
      entries_pte_U[entries_pte_U__T_17_addr] <= entries_pte_U__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_18_en & entries_pte_U__T_18_mask) begin
      entries_pte_U[entries_pte_U__T_18_addr] <= entries_pte_U__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_19_en & entries_pte_U__T_19_mask) begin
      entries_pte_U[entries_pte_U__T_19_addr] <= entries_pte_U__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_20_en & entries_pte_U__T_20_mask) begin
      entries_pte_U[entries_pte_U__T_20_addr] <= entries_pte_U__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_21_en & entries_pte_U__T_21_mask) begin
      entries_pte_U[entries_pte_U__T_21_addr] <= entries_pte_U__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_22_en & entries_pte_U__T_22_mask) begin
      entries_pte_U[entries_pte_U__T_22_addr] <= entries_pte_U__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_23_en & entries_pte_U__T_23_mask) begin
      entries_pte_U[entries_pte_U__T_23_addr] <= entries_pte_U__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_24_en & entries_pte_U__T_24_mask) begin
      entries_pte_U[entries_pte_U__T_24_addr] <= entries_pte_U__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_25_en & entries_pte_U__T_25_mask) begin
      entries_pte_U[entries_pte_U__T_25_addr] <= entries_pte_U__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_26_en & entries_pte_U__T_26_mask) begin
      entries_pte_U[entries_pte_U__T_26_addr] <= entries_pte_U__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_27_en & entries_pte_U__T_27_mask) begin
      entries_pte_U[entries_pte_U__T_27_addr] <= entries_pte_U__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_28_en & entries_pte_U__T_28_mask) begin
      entries_pte_U[entries_pte_U__T_28_addr] <= entries_pte_U__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_29_en & entries_pte_U__T_29_mask) begin
      entries_pte_U[entries_pte_U__T_29_addr] <= entries_pte_U__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_30_en & entries_pte_U__T_30_mask) begin
      entries_pte_U[entries_pte_U__T_30_addr] <= entries_pte_U__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_31_en & entries_pte_U__T_31_mask) begin
      entries_pte_U[entries_pte_U__T_31_addr] <= entries_pte_U__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_32_en & entries_pte_U__T_32_mask) begin
      entries_pte_U[entries_pte_U__T_32_addr] <= entries_pte_U__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_33_en & entries_pte_U__T_33_mask) begin
      entries_pte_U[entries_pte_U__T_33_addr] <= entries_pte_U__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_34_en & entries_pte_U__T_34_mask) begin
      entries_pte_U[entries_pte_U__T_34_addr] <= entries_pte_U__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_57_en & entries_pte_U__T_57_mask) begin
      entries_pte_U[entries_pte_U__T_57_addr] <= entries_pte_U__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_58_en & entries_pte_U__T_58_mask) begin
      entries_pte_U[entries_pte_U__T_58_addr] <= entries_pte_U__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_59_en & entries_pte_U__T_59_mask) begin
      entries_pte_U[entries_pte_U__T_59_addr] <= entries_pte_U__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_U__T_65_en & entries_pte_U__T_65_mask) begin
      entries_pte_U[entries_pte_U__T_65_addr] <= entries_pte_U__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_3_en & entries_pte_X__T_3_mask) begin
      entries_pte_X[entries_pte_X__T_3_addr] <= entries_pte_X__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_4_en & entries_pte_X__T_4_mask) begin
      entries_pte_X[entries_pte_X__T_4_addr] <= entries_pte_X__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_5_en & entries_pte_X__T_5_mask) begin
      entries_pte_X[entries_pte_X__T_5_addr] <= entries_pte_X__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_6_en & entries_pte_X__T_6_mask) begin
      entries_pte_X[entries_pte_X__T_6_addr] <= entries_pte_X__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_7_en & entries_pte_X__T_7_mask) begin
      entries_pte_X[entries_pte_X__T_7_addr] <= entries_pte_X__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_8_en & entries_pte_X__T_8_mask) begin
      entries_pte_X[entries_pte_X__T_8_addr] <= entries_pte_X__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_9_en & entries_pte_X__T_9_mask) begin
      entries_pte_X[entries_pte_X__T_9_addr] <= entries_pte_X__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_10_en & entries_pte_X__T_10_mask) begin
      entries_pte_X[entries_pte_X__T_10_addr] <= entries_pte_X__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_11_en & entries_pte_X__T_11_mask) begin
      entries_pte_X[entries_pte_X__T_11_addr] <= entries_pte_X__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_12_en & entries_pte_X__T_12_mask) begin
      entries_pte_X[entries_pte_X__T_12_addr] <= entries_pte_X__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_13_en & entries_pte_X__T_13_mask) begin
      entries_pte_X[entries_pte_X__T_13_addr] <= entries_pte_X__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_14_en & entries_pte_X__T_14_mask) begin
      entries_pte_X[entries_pte_X__T_14_addr] <= entries_pte_X__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_15_en & entries_pte_X__T_15_mask) begin
      entries_pte_X[entries_pte_X__T_15_addr] <= entries_pte_X__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_16_en & entries_pte_X__T_16_mask) begin
      entries_pte_X[entries_pte_X__T_16_addr] <= entries_pte_X__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_17_en & entries_pte_X__T_17_mask) begin
      entries_pte_X[entries_pte_X__T_17_addr] <= entries_pte_X__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_18_en & entries_pte_X__T_18_mask) begin
      entries_pte_X[entries_pte_X__T_18_addr] <= entries_pte_X__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_19_en & entries_pte_X__T_19_mask) begin
      entries_pte_X[entries_pte_X__T_19_addr] <= entries_pte_X__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_20_en & entries_pte_X__T_20_mask) begin
      entries_pte_X[entries_pte_X__T_20_addr] <= entries_pte_X__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_21_en & entries_pte_X__T_21_mask) begin
      entries_pte_X[entries_pte_X__T_21_addr] <= entries_pte_X__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_22_en & entries_pte_X__T_22_mask) begin
      entries_pte_X[entries_pte_X__T_22_addr] <= entries_pte_X__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_23_en & entries_pte_X__T_23_mask) begin
      entries_pte_X[entries_pte_X__T_23_addr] <= entries_pte_X__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_24_en & entries_pte_X__T_24_mask) begin
      entries_pte_X[entries_pte_X__T_24_addr] <= entries_pte_X__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_25_en & entries_pte_X__T_25_mask) begin
      entries_pte_X[entries_pte_X__T_25_addr] <= entries_pte_X__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_26_en & entries_pte_X__T_26_mask) begin
      entries_pte_X[entries_pte_X__T_26_addr] <= entries_pte_X__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_27_en & entries_pte_X__T_27_mask) begin
      entries_pte_X[entries_pte_X__T_27_addr] <= entries_pte_X__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_28_en & entries_pte_X__T_28_mask) begin
      entries_pte_X[entries_pte_X__T_28_addr] <= entries_pte_X__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_29_en & entries_pte_X__T_29_mask) begin
      entries_pte_X[entries_pte_X__T_29_addr] <= entries_pte_X__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_30_en & entries_pte_X__T_30_mask) begin
      entries_pte_X[entries_pte_X__T_30_addr] <= entries_pte_X__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_31_en & entries_pte_X__T_31_mask) begin
      entries_pte_X[entries_pte_X__T_31_addr] <= entries_pte_X__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_32_en & entries_pte_X__T_32_mask) begin
      entries_pte_X[entries_pte_X__T_32_addr] <= entries_pte_X__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_33_en & entries_pte_X__T_33_mask) begin
      entries_pte_X[entries_pte_X__T_33_addr] <= entries_pte_X__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_34_en & entries_pte_X__T_34_mask) begin
      entries_pte_X[entries_pte_X__T_34_addr] <= entries_pte_X__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_57_en & entries_pte_X__T_57_mask) begin
      entries_pte_X[entries_pte_X__T_57_addr] <= entries_pte_X__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_58_en & entries_pte_X__T_58_mask) begin
      entries_pte_X[entries_pte_X__T_58_addr] <= entries_pte_X__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_59_en & entries_pte_X__T_59_mask) begin
      entries_pte_X[entries_pte_X__T_59_addr] <= entries_pte_X__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_X__T_65_en & entries_pte_X__T_65_mask) begin
      entries_pte_X[entries_pte_X__T_65_addr] <= entries_pte_X__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_3_en & entries_pte_W__T_3_mask) begin
      entries_pte_W[entries_pte_W__T_3_addr] <= entries_pte_W__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_4_en & entries_pte_W__T_4_mask) begin
      entries_pte_W[entries_pte_W__T_4_addr] <= entries_pte_W__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_5_en & entries_pte_W__T_5_mask) begin
      entries_pte_W[entries_pte_W__T_5_addr] <= entries_pte_W__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_6_en & entries_pte_W__T_6_mask) begin
      entries_pte_W[entries_pte_W__T_6_addr] <= entries_pte_W__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_7_en & entries_pte_W__T_7_mask) begin
      entries_pte_W[entries_pte_W__T_7_addr] <= entries_pte_W__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_8_en & entries_pte_W__T_8_mask) begin
      entries_pte_W[entries_pte_W__T_8_addr] <= entries_pte_W__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_9_en & entries_pte_W__T_9_mask) begin
      entries_pte_W[entries_pte_W__T_9_addr] <= entries_pte_W__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_10_en & entries_pte_W__T_10_mask) begin
      entries_pte_W[entries_pte_W__T_10_addr] <= entries_pte_W__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_11_en & entries_pte_W__T_11_mask) begin
      entries_pte_W[entries_pte_W__T_11_addr] <= entries_pte_W__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_12_en & entries_pte_W__T_12_mask) begin
      entries_pte_W[entries_pte_W__T_12_addr] <= entries_pte_W__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_13_en & entries_pte_W__T_13_mask) begin
      entries_pte_W[entries_pte_W__T_13_addr] <= entries_pte_W__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_14_en & entries_pte_W__T_14_mask) begin
      entries_pte_W[entries_pte_W__T_14_addr] <= entries_pte_W__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_15_en & entries_pte_W__T_15_mask) begin
      entries_pte_W[entries_pte_W__T_15_addr] <= entries_pte_W__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_16_en & entries_pte_W__T_16_mask) begin
      entries_pte_W[entries_pte_W__T_16_addr] <= entries_pte_W__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_17_en & entries_pte_W__T_17_mask) begin
      entries_pte_W[entries_pte_W__T_17_addr] <= entries_pte_W__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_18_en & entries_pte_W__T_18_mask) begin
      entries_pte_W[entries_pte_W__T_18_addr] <= entries_pte_W__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_19_en & entries_pte_W__T_19_mask) begin
      entries_pte_W[entries_pte_W__T_19_addr] <= entries_pte_W__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_20_en & entries_pte_W__T_20_mask) begin
      entries_pte_W[entries_pte_W__T_20_addr] <= entries_pte_W__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_21_en & entries_pte_W__T_21_mask) begin
      entries_pte_W[entries_pte_W__T_21_addr] <= entries_pte_W__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_22_en & entries_pte_W__T_22_mask) begin
      entries_pte_W[entries_pte_W__T_22_addr] <= entries_pte_W__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_23_en & entries_pte_W__T_23_mask) begin
      entries_pte_W[entries_pte_W__T_23_addr] <= entries_pte_W__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_24_en & entries_pte_W__T_24_mask) begin
      entries_pte_W[entries_pte_W__T_24_addr] <= entries_pte_W__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_25_en & entries_pte_W__T_25_mask) begin
      entries_pte_W[entries_pte_W__T_25_addr] <= entries_pte_W__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_26_en & entries_pte_W__T_26_mask) begin
      entries_pte_W[entries_pte_W__T_26_addr] <= entries_pte_W__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_27_en & entries_pte_W__T_27_mask) begin
      entries_pte_W[entries_pte_W__T_27_addr] <= entries_pte_W__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_28_en & entries_pte_W__T_28_mask) begin
      entries_pte_W[entries_pte_W__T_28_addr] <= entries_pte_W__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_29_en & entries_pte_W__T_29_mask) begin
      entries_pte_W[entries_pte_W__T_29_addr] <= entries_pte_W__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_30_en & entries_pte_W__T_30_mask) begin
      entries_pte_W[entries_pte_W__T_30_addr] <= entries_pte_W__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_31_en & entries_pte_W__T_31_mask) begin
      entries_pte_W[entries_pte_W__T_31_addr] <= entries_pte_W__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_32_en & entries_pte_W__T_32_mask) begin
      entries_pte_W[entries_pte_W__T_32_addr] <= entries_pte_W__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_33_en & entries_pte_W__T_33_mask) begin
      entries_pte_W[entries_pte_W__T_33_addr] <= entries_pte_W__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_34_en & entries_pte_W__T_34_mask) begin
      entries_pte_W[entries_pte_W__T_34_addr] <= entries_pte_W__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_57_en & entries_pte_W__T_57_mask) begin
      entries_pte_W[entries_pte_W__T_57_addr] <= entries_pte_W__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_58_en & entries_pte_W__T_58_mask) begin
      entries_pte_W[entries_pte_W__T_58_addr] <= entries_pte_W__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_59_en & entries_pte_W__T_59_mask) begin
      entries_pte_W[entries_pte_W__T_59_addr] <= entries_pte_W__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_W__T_65_en & entries_pte_W__T_65_mask) begin
      entries_pte_W[entries_pte_W__T_65_addr] <= entries_pte_W__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_3_en & entries_pte_R__T_3_mask) begin
      entries_pte_R[entries_pte_R__T_3_addr] <= entries_pte_R__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_4_en & entries_pte_R__T_4_mask) begin
      entries_pte_R[entries_pte_R__T_4_addr] <= entries_pte_R__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_5_en & entries_pte_R__T_5_mask) begin
      entries_pte_R[entries_pte_R__T_5_addr] <= entries_pte_R__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_6_en & entries_pte_R__T_6_mask) begin
      entries_pte_R[entries_pte_R__T_6_addr] <= entries_pte_R__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_7_en & entries_pte_R__T_7_mask) begin
      entries_pte_R[entries_pte_R__T_7_addr] <= entries_pte_R__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_8_en & entries_pte_R__T_8_mask) begin
      entries_pte_R[entries_pte_R__T_8_addr] <= entries_pte_R__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_9_en & entries_pte_R__T_9_mask) begin
      entries_pte_R[entries_pte_R__T_9_addr] <= entries_pte_R__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_10_en & entries_pte_R__T_10_mask) begin
      entries_pte_R[entries_pte_R__T_10_addr] <= entries_pte_R__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_11_en & entries_pte_R__T_11_mask) begin
      entries_pte_R[entries_pte_R__T_11_addr] <= entries_pte_R__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_12_en & entries_pte_R__T_12_mask) begin
      entries_pte_R[entries_pte_R__T_12_addr] <= entries_pte_R__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_13_en & entries_pte_R__T_13_mask) begin
      entries_pte_R[entries_pte_R__T_13_addr] <= entries_pte_R__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_14_en & entries_pte_R__T_14_mask) begin
      entries_pte_R[entries_pte_R__T_14_addr] <= entries_pte_R__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_15_en & entries_pte_R__T_15_mask) begin
      entries_pte_R[entries_pte_R__T_15_addr] <= entries_pte_R__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_16_en & entries_pte_R__T_16_mask) begin
      entries_pte_R[entries_pte_R__T_16_addr] <= entries_pte_R__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_17_en & entries_pte_R__T_17_mask) begin
      entries_pte_R[entries_pte_R__T_17_addr] <= entries_pte_R__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_18_en & entries_pte_R__T_18_mask) begin
      entries_pte_R[entries_pte_R__T_18_addr] <= entries_pte_R__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_19_en & entries_pte_R__T_19_mask) begin
      entries_pte_R[entries_pte_R__T_19_addr] <= entries_pte_R__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_20_en & entries_pte_R__T_20_mask) begin
      entries_pte_R[entries_pte_R__T_20_addr] <= entries_pte_R__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_21_en & entries_pte_R__T_21_mask) begin
      entries_pte_R[entries_pte_R__T_21_addr] <= entries_pte_R__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_22_en & entries_pte_R__T_22_mask) begin
      entries_pte_R[entries_pte_R__T_22_addr] <= entries_pte_R__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_23_en & entries_pte_R__T_23_mask) begin
      entries_pte_R[entries_pte_R__T_23_addr] <= entries_pte_R__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_24_en & entries_pte_R__T_24_mask) begin
      entries_pte_R[entries_pte_R__T_24_addr] <= entries_pte_R__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_25_en & entries_pte_R__T_25_mask) begin
      entries_pte_R[entries_pte_R__T_25_addr] <= entries_pte_R__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_26_en & entries_pte_R__T_26_mask) begin
      entries_pte_R[entries_pte_R__T_26_addr] <= entries_pte_R__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_27_en & entries_pte_R__T_27_mask) begin
      entries_pte_R[entries_pte_R__T_27_addr] <= entries_pte_R__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_28_en & entries_pte_R__T_28_mask) begin
      entries_pte_R[entries_pte_R__T_28_addr] <= entries_pte_R__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_29_en & entries_pte_R__T_29_mask) begin
      entries_pte_R[entries_pte_R__T_29_addr] <= entries_pte_R__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_30_en & entries_pte_R__T_30_mask) begin
      entries_pte_R[entries_pte_R__T_30_addr] <= entries_pte_R__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_31_en & entries_pte_R__T_31_mask) begin
      entries_pte_R[entries_pte_R__T_31_addr] <= entries_pte_R__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_32_en & entries_pte_R__T_32_mask) begin
      entries_pte_R[entries_pte_R__T_32_addr] <= entries_pte_R__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_33_en & entries_pte_R__T_33_mask) begin
      entries_pte_R[entries_pte_R__T_33_addr] <= entries_pte_R__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_34_en & entries_pte_R__T_34_mask) begin
      entries_pte_R[entries_pte_R__T_34_addr] <= entries_pte_R__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_57_en & entries_pte_R__T_57_mask) begin
      entries_pte_R[entries_pte_R__T_57_addr] <= entries_pte_R__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_58_en & entries_pte_R__T_58_mask) begin
      entries_pte_R[entries_pte_R__T_58_addr] <= entries_pte_R__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_59_en & entries_pte_R__T_59_mask) begin
      entries_pte_R[entries_pte_R__T_59_addr] <= entries_pte_R__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_R__T_65_en & entries_pte_R__T_65_mask) begin
      entries_pte_R[entries_pte_R__T_65_addr] <= entries_pte_R__T_65_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_3_en & entries_pte_V__T_3_mask) begin
      entries_pte_V[entries_pte_V__T_3_addr] <= entries_pte_V__T_3_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_4_en & entries_pte_V__T_4_mask) begin
      entries_pte_V[entries_pte_V__T_4_addr] <= entries_pte_V__T_4_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_5_en & entries_pte_V__T_5_mask) begin
      entries_pte_V[entries_pte_V__T_5_addr] <= entries_pte_V__T_5_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_6_en & entries_pte_V__T_6_mask) begin
      entries_pte_V[entries_pte_V__T_6_addr] <= entries_pte_V__T_6_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_7_en & entries_pte_V__T_7_mask) begin
      entries_pte_V[entries_pte_V__T_7_addr] <= entries_pte_V__T_7_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_8_en & entries_pte_V__T_8_mask) begin
      entries_pte_V[entries_pte_V__T_8_addr] <= entries_pte_V__T_8_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_9_en & entries_pte_V__T_9_mask) begin
      entries_pte_V[entries_pte_V__T_9_addr] <= entries_pte_V__T_9_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_10_en & entries_pte_V__T_10_mask) begin
      entries_pte_V[entries_pte_V__T_10_addr] <= entries_pte_V__T_10_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_11_en & entries_pte_V__T_11_mask) begin
      entries_pte_V[entries_pte_V__T_11_addr] <= entries_pte_V__T_11_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_12_en & entries_pte_V__T_12_mask) begin
      entries_pte_V[entries_pte_V__T_12_addr] <= entries_pte_V__T_12_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_13_en & entries_pte_V__T_13_mask) begin
      entries_pte_V[entries_pte_V__T_13_addr] <= entries_pte_V__T_13_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_14_en & entries_pte_V__T_14_mask) begin
      entries_pte_V[entries_pte_V__T_14_addr] <= entries_pte_V__T_14_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_15_en & entries_pte_V__T_15_mask) begin
      entries_pte_V[entries_pte_V__T_15_addr] <= entries_pte_V__T_15_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_16_en & entries_pte_V__T_16_mask) begin
      entries_pte_V[entries_pte_V__T_16_addr] <= entries_pte_V__T_16_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_17_en & entries_pte_V__T_17_mask) begin
      entries_pte_V[entries_pte_V__T_17_addr] <= entries_pte_V__T_17_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_18_en & entries_pte_V__T_18_mask) begin
      entries_pte_V[entries_pte_V__T_18_addr] <= entries_pte_V__T_18_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_19_en & entries_pte_V__T_19_mask) begin
      entries_pte_V[entries_pte_V__T_19_addr] <= entries_pte_V__T_19_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_20_en & entries_pte_V__T_20_mask) begin
      entries_pte_V[entries_pte_V__T_20_addr] <= entries_pte_V__T_20_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_21_en & entries_pte_V__T_21_mask) begin
      entries_pte_V[entries_pte_V__T_21_addr] <= entries_pte_V__T_21_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_22_en & entries_pte_V__T_22_mask) begin
      entries_pte_V[entries_pte_V__T_22_addr] <= entries_pte_V__T_22_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_23_en & entries_pte_V__T_23_mask) begin
      entries_pte_V[entries_pte_V__T_23_addr] <= entries_pte_V__T_23_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_24_en & entries_pte_V__T_24_mask) begin
      entries_pte_V[entries_pte_V__T_24_addr] <= entries_pte_V__T_24_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_25_en & entries_pte_V__T_25_mask) begin
      entries_pte_V[entries_pte_V__T_25_addr] <= entries_pte_V__T_25_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_26_en & entries_pte_V__T_26_mask) begin
      entries_pte_V[entries_pte_V__T_26_addr] <= entries_pte_V__T_26_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_27_en & entries_pte_V__T_27_mask) begin
      entries_pte_V[entries_pte_V__T_27_addr] <= entries_pte_V__T_27_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_28_en & entries_pte_V__T_28_mask) begin
      entries_pte_V[entries_pte_V__T_28_addr] <= entries_pte_V__T_28_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_29_en & entries_pte_V__T_29_mask) begin
      entries_pte_V[entries_pte_V__T_29_addr] <= entries_pte_V__T_29_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_30_en & entries_pte_V__T_30_mask) begin
      entries_pte_V[entries_pte_V__T_30_addr] <= entries_pte_V__T_30_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_31_en & entries_pte_V__T_31_mask) begin
      entries_pte_V[entries_pte_V__T_31_addr] <= entries_pte_V__T_31_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_32_en & entries_pte_V__T_32_mask) begin
      entries_pte_V[entries_pte_V__T_32_addr] <= entries_pte_V__T_32_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_33_en & entries_pte_V__T_33_mask) begin
      entries_pte_V[entries_pte_V__T_33_addr] <= entries_pte_V__T_33_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_34_en & entries_pte_V__T_34_mask) begin
      entries_pte_V[entries_pte_V__T_34_addr] <= entries_pte_V__T_34_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_57_en & entries_pte_V__T_57_mask) begin
      entries_pte_V[entries_pte_V__T_57_addr] <= entries_pte_V__T_57_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_58_en & entries_pte_V__T_58_mask) begin
      entries_pte_V[entries_pte_V__T_58_addr] <= entries_pte_V__T_58_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_59_en & entries_pte_V__T_59_mask) begin
      entries_pte_V[entries_pte_V__T_59_addr] <= entries_pte_V__T_59_data; // @[TLB.scala 38:20]
    end
    if(entries_pte_V__T_65_en & entries_pte_V__T_65_mask) begin
      entries_pte_V[entries_pte_V__T_65_addr] <= entries_pte_V__T_65_data; // @[TLB.scala 38:20]
    end
  end
endmodule
module MMU(
  input         clock,
  input         reset,
  input  [31:0] io_iff_addr,
  input  [3:0]  io_iff_mode,
  output [31:0] io_iff_rdata,
  output        io_iff_ok,
  output        io_iff_pageFault,
  input  [31:0] io_mem_addr,
  input  [3:0]  io_mem_mode,
  input  [31:0] io_mem_wdata,
  output [31:0] io_mem_rdata,
  output        io_mem_ok,
  output        io_mem_pageFault,
  input  [31:0] io_csr_satp,
  input         io_csr_flush_one,
  input         io_csr_flush_all,
  input  [31:0] io_csr_flush_addr,
  input  [1:0]  io_csr_priv,
  input         io_csr_mxr,
  input         io_csr_sum,
  output [31:0] io_dev_if__addr,
  output [3:0]  io_dev_if__mode,
  input  [31:0] io_dev_if__rdata,
  input         io_dev_if__ok,
  output [31:0] io_dev_mem_addr,
  output [3:0]  io_dev_mem_mode,
  output [31:0] io_dev_mem_wdata,
  input  [31:0] io_dev_mem_rdata,
  input         io_dev_mem_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  ptw_clock; // @[MMU.scala 17:19]
  wire  ptw_reset; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_root_p2; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_root_p1; // @[MMU.scala 17:19]
  wire  ptw_io_req_ready; // @[MMU.scala 17:19]
  wire  ptw_io_req_valid; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_req_bits_p2; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_req_bits_p1; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_ready; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_valid; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_rsp_bits_ppn_p2; // @[MMU.scala 17:19]
  wire [9:0] ptw_io_rsp_bits_ppn_p1; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_bits_U; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_bits_X; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_bits_W; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_bits_R; // @[MMU.scala 17:19]
  wire  ptw_io_rsp_bits_V; // @[MMU.scala 17:19]
  wire [31:0] ptw_io_mem_addr; // @[MMU.scala 17:19]
  wire [3:0] ptw_io_mem_mode; // @[MMU.scala 17:19]
  wire [31:0] ptw_io_mem_rdata; // @[MMU.scala 17:19]
  wire  ptw_io_mem_ok; // @[MMU.scala 17:19]
  wire  tlb_clock; // @[MMU.scala 18:19]
  wire  tlb_reset; // @[MMU.scala 18:19]
  wire  tlb_io_query_req_valid; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query_req_bits_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query_req_bits_p1; // @[MMU.scala 18:19]
  wire  tlb_io_query_rsp_valid; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query_rsp_bits_ppn_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query_rsp_bits_ppn_p1; // @[MMU.scala 18:19]
  wire  tlb_io_query_rsp_bits_U; // @[MMU.scala 18:19]
  wire  tlb_io_query_rsp_bits_X; // @[MMU.scala 18:19]
  wire  tlb_io_query_rsp_bits_V; // @[MMU.scala 18:19]
  wire  tlb_io_query2_req_valid; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query2_req_bits_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query2_req_bits_p1; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_valid; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query2_rsp_bits_ppn_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_query2_rsp_bits_ppn_p1; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_bits_U; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_bits_X; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_bits_W; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_bits_R; // @[MMU.scala 18:19]
  wire  tlb_io_query2_rsp_bits_V; // @[MMU.scala 18:19]
  wire [1:0] tlb_io_modify_mode; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_modify_vpn_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_modify_vpn_p1; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_modify_pte_ppn_p2; // @[MMU.scala 18:19]
  wire [9:0] tlb_io_modify_pte_ppn_p1; // @[MMU.scala 18:19]
  wire  tlb_io_modify_pte_U; // @[MMU.scala 18:19]
  wire  tlb_io_modify_pte_X; // @[MMU.scala 18:19]
  wire  tlb_io_modify_pte_W; // @[MMU.scala 18:19]
  wire  tlb_io_modify_pte_R; // @[MMU.scala 18:19]
  wire  tlb_io_modify_pte_V; // @[MMU.scala 18:19]
  wire  _T = io_iff_mode == 4'h0; // @[Bundles.scala 57:20]
  wire  _T_1 = _T | io_iff_ok; // @[Bundles.scala 57:36]
  wire  _T_2 = io_mem_mode == 4'h0; // @[Bundles.scala 57:20]
  wire  _T_3 = _T_2 | io_mem_ok; // @[Bundles.scala 57:36]
  wire  ready = _T_1 & _T_3; // @[MMU.scala 22:28]
  reg [31:0] csr_satp; // @[MMU.scala 24:20]
  reg [1:0] csr_priv; // @[MMU.scala 24:20]
  reg  csr_mxr; // @[MMU.scala 24:20]
  reg  csr_sum; // @[MMU.scala 24:20]
  reg  log_flush_one; // @[MMU.scala 32:26]
  reg  log_flush_all; // @[MMU.scala 32:26]
  reg [31:0] log_flush_addr; // @[MMU.scala 32:26]
  wire  _T_6 = io_csr_flush_one | io_csr_flush_all; // @[Bundles.scala 68:19]
  wire [31:0] _GEN_7 = _T_6 ? io_csr_flush_addr : log_flush_addr; // @[MMU.scala 33:28]
  wire  _GEN_8 = _T_6 ? io_csr_flush_all : log_flush_all; // @[MMU.scala 33:28]
  wire  _GEN_9 = _T_6 ? io_csr_flush_one : log_flush_one; // @[MMU.scala 33:28]
  wire  _T_9 = csr_priv != 2'h3; // @[MMU.scala 40:41]
  wire  enable = csr_satp[31] & _T_9; // @[MMU.scala 40:29]
  wire  _T_16 = io_iff_mode != 4'h0; // @[MMU.scala 50:31]
  wire [31:0] _T_25 = {tlb_io_query_rsp_bits_ppn_p2,tlb_io_query_rsp_bits_ppn_p1,io_iff_addr[11:0]}; // @[PTW.scala 12:53]
  wire  _T_26 = io_dev_if__ok & tlb_io_query_rsp_valid; // @[MMU.scala 57:22]
  wire  _T_27 = ~tlb_io_query_rsp_valid; // @[TLB.scala 9:27]
  wire  _T_28 = tlb_io_query_req_valid & _T_27; // @[TLB.scala 9:24]
  wire [3:0] _GEN_10 = io_iff_pageFault ? 4'h0 : io_iff_mode; // @[MMU.scala 63:31]
  wire [31:0] _GEN_12 = io_iff_pageFault ? 32'h0 : _T_25; // @[MMU.scala 63:31]
  wire  _GEN_13 = io_iff_pageFault | _T_26; // @[MMU.scala 63:31]
  wire [3:0] _GEN_14 = _T_28 ? 4'h0 : _GEN_10; // @[MMU.scala 60:20]
  wire  _GEN_15 = _T_28 ? 1'h0 : _GEN_13; // @[MMU.scala 60:20]
  wire [31:0] _GEN_17 = _T_28 ? _T_25 : _GEN_12; // @[MMU.scala 60:20]
  wire  _T_29 = io_mem_mode != 4'h0; // @[MMU.scala 50:31]
  wire [31:0] _T_37 = {tlb_io_query2_rsp_bits_ppn_p2,tlb_io_query2_rsp_bits_ppn_p1,io_mem_addr[11:0]}; // @[PTW.scala 12:53]
  wire  _T_38 = io_dev_mem_ok & tlb_io_query2_rsp_valid; // @[MMU.scala 57:22]
  wire  _T_39 = ~tlb_io_query2_rsp_valid; // @[TLB.scala 9:27]
  wire  _T_40 = tlb_io_query2_req_valid & _T_39; // @[TLB.scala 9:24]
  wire [3:0] _GEN_18 = io_mem_pageFault ? 4'h0 : io_mem_mode; // @[MMU.scala 63:31]
  wire [31:0] _GEN_19 = io_mem_pageFault ? 32'h0 : io_mem_wdata; // @[MMU.scala 63:31]
  wire [31:0] _GEN_20 = io_mem_pageFault ? 32'h0 : _T_37; // @[MMU.scala 63:31]
  wire  _GEN_21 = io_mem_pageFault | _T_38; // @[MMU.scala 63:31]
  wire [3:0] _GEN_22 = _T_40 ? 4'h0 : _GEN_18; // @[MMU.scala 60:20]
  wire  _GEN_23 = _T_40 ? 1'h0 : _GEN_21; // @[MMU.scala 60:20]
  wire  _T_41 = tlb_io_query_rsp_bits_V & tlb_io_query_rsp_bits_X; // @[MMU.scala 76:31]
  wire  _T_42 = ~_T_41; // @[MMU.scala 76:18]
  wire  _T_43 = csr_priv == 2'h0; // @[MMU.scala 77:27]
  wire  _T_44 = ~tlb_io_query_rsp_bits_U; // @[MMU.scala 77:41]
  wire  _T_45 = _T_43 & _T_44; // @[MMU.scala 77:38]
  wire  _T_46 = enable & tlb_io_query_rsp_valid; // @[MMU.scala 78:32]
  wire  _T_48 = _T_46 & _T_16; // @[MMU.scala 78:45]
  wire  _T_49 = _T_42 | _T_45; // @[MMU.scala 78:87]
  wire  _T_52 = ~io_mem_mode[3]; // @[Const.scala 23:32]
  wire  _T_53 = |io_mem_mode; // @[Const.scala 23:43]
  wire  _T_54 = _T_52 & _T_53; // @[Const.scala 23:38]
  wire  _T_55 = tlb_io_query2_rsp_bits_X & csr_mxr; // @[MMU.scala 82:92]
  wire  _T_56 = tlb_io_query2_rsp_bits_R | _T_55; // @[MMU.scala 82:78]
  wire  _T_57 = tlb_io_query2_rsp_bits_V & _T_56; // @[MMU.scala 82:63]
  wire  _T_58 = ~_T_57; // @[MMU.scala 82:50]
  wire  _T_59 = _T_54 & _T_58; // @[MMU.scala 82:47]
  wire  _T_61 = tlb_io_query2_rsp_bits_V & tlb_io_query2_rsp_bits_W; // @[MMU.scala 83:64]
  wire  _T_62 = ~_T_61; // @[MMU.scala 83:51]
  wire  _T_63 = io_mem_mode[3] & _T_62; // @[MMU.scala 83:48]
  wire  _T_65 = ~tlb_io_query2_rsp_bits_U; // @[MMU.scala 84:42]
  wire  _T_66 = _T_43 & _T_65; // @[MMU.scala 84:39]
  wire  _T_67 = csr_priv == 2'h1; // @[MMU.scala 85:28]
  wire  _T_68 = ~csr_sum; // @[MMU.scala 85:42]
  wire  _T_69 = _T_67 & _T_68; // @[MMU.scala 85:39]
  wire  _T_70 = _T_69 & tlb_io_query2_rsp_bits_U; // @[MMU.scala 85:51]
  wire  _T_71 = enable & tlb_io_query2_rsp_valid; // @[MMU.scala 86:32]
  wire  _T_73 = _T_71 & _T_29; // @[MMU.scala 86:45]
  wire  _T_74 = _T_59 | _T_63; // @[MMU.scala 86:87]
  wire  _T_75 = _T_74 | _T_66; // @[MMU.scala 86:98]
  wire  _T_76 = _T_75 | _T_70; // @[MMU.scala 86:108]
  reg  status; // @[MMU.scala 100:23]
  reg [9:0] ptw_vpn_p2; // @[MMU.scala 101:24]
  reg [9:0] ptw_vpn_p1; // @[MMU.scala 101:24]
  wire  _T_81 = ~status; // @[Conditional.scala 37:30]
  wire  _T_82 = io_dev_mem_mode == 4'h0; // @[Bundles.scala 57:20]
  wire  _T_83 = _T_82 | io_dev_mem_ok; // @[Bundles.scala 57:36]
  wire  _T_86 = _T_28 & _T_83; // @[MMU.scala 112:23]
  wire  _T_87 = _T_86 & ptw_io_req_ready; // @[MMU.scala 112:37]
  wire [9:0] _GEN_27 = _T_87 ? tlb_io_query_req_bits_p1 : 10'h0; // @[MMU.scala 112:58]
  wire [9:0] _GEN_28 = _T_87 ? tlb_io_query_req_bits_p2 : 10'h0; // @[MMU.scala 112:58]
  wire  _GEN_29 = _T_87 | status; // @[MMU.scala 112:58]
  wire  _T_88 = io_dev_if__mode == 4'h0; // @[Bundles.scala 57:20]
  wire  _T_89 = _T_88 | io_dev_if__ok; // @[Bundles.scala 57:36]
  wire  _T_92 = _T_40 & _T_89; // @[MMU.scala 112:23]
  wire  _T_93 = _T_92 & ptw_io_req_ready; // @[MMU.scala 112:37]
  wire  _GEN_32 = _T_93 | _T_87; // @[MMU.scala 112:58]
  wire [9:0] _GEN_33 = _T_93 ? tlb_io_query2_req_bits_p1 : _GEN_27; // @[MMU.scala 112:58]
  wire [9:0] _GEN_34 = _T_93 ? tlb_io_query2_req_bits_p2 : _GEN_28; // @[MMU.scala 112:58]
  wire  _GEN_35 = _T_93 | _GEN_29; // @[MMU.scala 112:58]
  wire [1:0] _GEN_38 = _GEN_8 ? 2'h3 : 2'h0; // @[MMU.scala 127:31]
  wire [1:0] _GEN_39 = _GEN_9 ? 2'h2 : _GEN_38; // @[MMU.scala 124:25]
  wire [9:0] _GEN_40 = _GEN_9 ? _GEN_7[21:12] : 10'h0; // @[MMU.scala 124:25]
  wire [9:0] _GEN_41 = _GEN_9 ? _GEN_7[31:22] : 10'h0; // @[MMU.scala 124:25]
  wire [1:0] _GEN_42 = ready ? _GEN_39 : 2'h0; // @[MMU.scala 123:19]
  wire [9:0] _GEN_43 = ready ? _GEN_40 : 10'h0; // @[MMU.scala 123:19]
  wire [9:0] _GEN_44 = ready ? _GEN_41 : 10'h0; // @[MMU.scala 123:19]
  reg [31:0] _T_101; // @[MMU.scala 137:33]
  reg [3:0] _T_102; // @[MMU.scala 138:33]
  wire [1:0] _GEN_48 = ptw_io_rsp_valid ? 2'h1 : 2'h0; // @[MMU.scala 147:30]
  wire [9:0] _GEN_49 = ptw_io_rsp_valid ? ptw_vpn_p1 : 10'h0; // @[MMU.scala 147:30]
  wire [9:0] _GEN_50 = ptw_io_rsp_valid ? ptw_vpn_p2 : 10'h0; // @[MMU.scala 147:30]
  wire  _GEN_51 = ptw_io_rsp_valid & ptw_io_rsp_bits_V; // @[MMU.scala 147:30]
  wire  _GEN_52 = ptw_io_rsp_valid & ptw_io_rsp_bits_R; // @[MMU.scala 147:30]
  wire  _GEN_53 = ptw_io_rsp_valid & ptw_io_rsp_bits_W; // @[MMU.scala 147:30]
  wire  _GEN_54 = ptw_io_rsp_valid & ptw_io_rsp_bits_X; // @[MMU.scala 147:30]
  wire  _GEN_55 = ptw_io_rsp_valid & ptw_io_rsp_bits_U; // @[MMU.scala 147:30]
  wire [9:0] _GEN_60 = ptw_io_rsp_valid ? ptw_io_rsp_bits_ppn_p1 : 10'h0; // @[MMU.scala 147:30]
  wire [9:0] _GEN_61 = ptw_io_rsp_valid ? ptw_io_rsp_bits_ppn_p2 : 10'h0; // @[MMU.scala 147:30]
  wire [31:0] _GEN_64 = status ? _T_101 : _GEN_17; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_65 = status ? _T_102 : _GEN_14; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_67 = status ? io_dev_if__rdata : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_68 = status & io_dev_if__ok; // @[Conditional.scala 39:67]
  wire  _GEN_69 = status ? 1'h0 : _GEN_15; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_70 = status ? 4'h0 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_71 = status ? 1'h0 : _GEN_23; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_73 = status ? _GEN_48 : 2'h0; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_74 = status ? _GEN_49 : 10'h0; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_75 = status ? _GEN_50 : 10'h0; // @[Conditional.scala 39:67]
  wire  _GEN_76 = status & _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_77 = status & _GEN_52; // @[Conditional.scala 39:67]
  wire  _GEN_78 = status & _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_79 = status & _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_80 = status & _GEN_55; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_85 = status ? _GEN_60 : 10'h0; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_86 = status ? _GEN_61 : 10'h0; // @[Conditional.scala 39:67]
  PTW ptw ( // @[MMU.scala 17:19]
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_root_p2(ptw_io_root_p2),
    .io_root_p1(ptw_io_root_p1),
    .io_req_ready(ptw_io_req_ready),
    .io_req_valid(ptw_io_req_valid),
    .io_req_bits_p2(ptw_io_req_bits_p2),
    .io_req_bits_p1(ptw_io_req_bits_p1),
    .io_rsp_ready(ptw_io_rsp_ready),
    .io_rsp_valid(ptw_io_rsp_valid),
    .io_rsp_bits_ppn_p2(ptw_io_rsp_bits_ppn_p2),
    .io_rsp_bits_ppn_p1(ptw_io_rsp_bits_ppn_p1),
    .io_rsp_bits_U(ptw_io_rsp_bits_U),
    .io_rsp_bits_X(ptw_io_rsp_bits_X),
    .io_rsp_bits_W(ptw_io_rsp_bits_W),
    .io_rsp_bits_R(ptw_io_rsp_bits_R),
    .io_rsp_bits_V(ptw_io_rsp_bits_V),
    .io_mem_addr(ptw_io_mem_addr),
    .io_mem_mode(ptw_io_mem_mode),
    .io_mem_rdata(ptw_io_mem_rdata),
    .io_mem_ok(ptw_io_mem_ok)
  );
  TLB tlb ( // @[MMU.scala 18:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_query_req_valid(tlb_io_query_req_valid),
    .io_query_req_bits_p2(tlb_io_query_req_bits_p2),
    .io_query_req_bits_p1(tlb_io_query_req_bits_p1),
    .io_query_rsp_valid(tlb_io_query_rsp_valid),
    .io_query_rsp_bits_ppn_p2(tlb_io_query_rsp_bits_ppn_p2),
    .io_query_rsp_bits_ppn_p1(tlb_io_query_rsp_bits_ppn_p1),
    .io_query_rsp_bits_U(tlb_io_query_rsp_bits_U),
    .io_query_rsp_bits_X(tlb_io_query_rsp_bits_X),
    .io_query_rsp_bits_V(tlb_io_query_rsp_bits_V),
    .io_query2_req_valid(tlb_io_query2_req_valid),
    .io_query2_req_bits_p2(tlb_io_query2_req_bits_p2),
    .io_query2_req_bits_p1(tlb_io_query2_req_bits_p1),
    .io_query2_rsp_valid(tlb_io_query2_rsp_valid),
    .io_query2_rsp_bits_ppn_p2(tlb_io_query2_rsp_bits_ppn_p2),
    .io_query2_rsp_bits_ppn_p1(tlb_io_query2_rsp_bits_ppn_p1),
    .io_query2_rsp_bits_U(tlb_io_query2_rsp_bits_U),
    .io_query2_rsp_bits_X(tlb_io_query2_rsp_bits_X),
    .io_query2_rsp_bits_W(tlb_io_query2_rsp_bits_W),
    .io_query2_rsp_bits_R(tlb_io_query2_rsp_bits_R),
    .io_query2_rsp_bits_V(tlb_io_query2_rsp_bits_V),
    .io_modify_mode(tlb_io_modify_mode),
    .io_modify_vpn_p2(tlb_io_modify_vpn_p2),
    .io_modify_vpn_p1(tlb_io_modify_vpn_p1),
    .io_modify_pte_ppn_p2(tlb_io_modify_pte_ppn_p2),
    .io_modify_pte_ppn_p1(tlb_io_modify_pte_ppn_p1),
    .io_modify_pte_U(tlb_io_modify_pte_U),
    .io_modify_pte_X(tlb_io_modify_pte_X),
    .io_modify_pte_W(tlb_io_modify_pte_W),
    .io_modify_pte_R(tlb_io_modify_pte_R),
    .io_modify_pte_V(tlb_io_modify_pte_V)
  );
  assign io_iff_rdata = io_dev_if__rdata; // @[MMU.scala 58:15]
  assign io_iff_ok = _T_81 ? _GEN_15 : _GEN_69; // @[MMU.scala 57:12 MMU.scala 62:14 MMU.scala 67:14 MMU.scala 143:17]
  assign io_iff_pageFault = _T_48 & _T_49; // @[MMU.scala 78:22]
  assign io_mem_rdata = io_dev_mem_rdata; // @[MMU.scala 58:15]
  assign io_mem_ok = _T_81 ? _GEN_23 : _GEN_71; // @[MMU.scala 57:12 MMU.scala 62:14 MMU.scala 67:14 MMU.scala 145:17]
  assign io_mem_pageFault = _T_73 & _T_76; // @[MMU.scala 86:22]
  assign io_dev_if__addr = _T_81 ? _GEN_17 : _GEN_64; // @[MMU.scala 55:14 MMU.scala 66:16 MMU.scala 137:23]
  assign io_dev_if__mode = _T_81 ? _GEN_14 : _GEN_65; // @[MMU.scala 53:14 MMU.scala 61:16 MMU.scala 64:16 MMU.scala 138:23]
  assign io_dev_mem_addr = _T_40 ? _T_37 : _GEN_20; // @[MMU.scala 55:14 MMU.scala 66:16]
  assign io_dev_mem_mode = _T_81 ? _GEN_22 : _GEN_70; // @[MMU.scala 53:14 MMU.scala 61:16 MMU.scala 64:16 MMU.scala 144:23]
  assign io_dev_mem_wdata = _T_40 ? io_mem_wdata : _GEN_19; // @[MMU.scala 54:15 MMU.scala 65:17]
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_root_p2 = csr_satp[19:10]; // @[MMU.scala 42:15]
  assign ptw_io_root_p1 = csr_satp[9:0]; // @[MMU.scala 42:15]
  assign ptw_io_req_valid = _T_81 & _GEN_32; // @[MMU.scala 104:20 MMU.scala 113:28 MMU.scala 113:28]
  assign ptw_io_req_bits_p2 = _T_81 ? _GEN_34 : 10'h0; // @[MMU.scala 105:19 MMU.scala 114:27 MMU.scala 114:27]
  assign ptw_io_req_bits_p1 = _T_81 ? _GEN_33 : 10'h0; // @[MMU.scala 105:19 MMU.scala 114:27 MMU.scala 114:27]
  assign ptw_io_rsp_ready = _T_81 ? 1'h0 : status; // @[MMU.scala 106:20 MMU.scala 146:24]
  assign ptw_io_mem_rdata = _T_81 ? 32'h0 : _GEN_67; // @[MMU.scala 45:14 MMU.scala 140:24]
  assign ptw_io_mem_ok = _T_81 ? 1'h0 : _GEN_68; // @[MMU.scala 45:14 MMU.scala 141:21]
  assign tlb_clock = clock;
  assign tlb_reset = ~enable; // @[MMU.scala 41:13]
  assign tlb_io_query_req_valid = io_iff_mode != 4'h0; // @[MMU.scala 50:19]
  assign tlb_io_query_req_bits_p2 = io_iff_addr[31:22]; // @[MMU.scala 51:18]
  assign tlb_io_query_req_bits_p1 = io_iff_addr[21:12]; // @[MMU.scala 51:18]
  assign tlb_io_query2_req_valid = io_mem_mode != 4'h0; // @[MMU.scala 50:19]
  assign tlb_io_query2_req_bits_p2 = io_mem_addr[31:22]; // @[MMU.scala 51:18]
  assign tlb_io_query2_req_bits_p1 = io_mem_addr[21:12]; // @[MMU.scala 51:18]
  assign tlb_io_modify_mode = _T_81 ? _GEN_42 : _GEN_73; // @[MMU.scala 107:17 MMU.scala 125:30 MMU.scala 128:30 MMU.scala 148:28]
  assign tlb_io_modify_vpn_p2 = _T_81 ? _GEN_44 : _GEN_75; // @[MMU.scala 107:17 MMU.scala 126:29 MMU.scala 149:27]
  assign tlb_io_modify_vpn_p1 = _T_81 ? _GEN_43 : _GEN_74; // @[MMU.scala 107:17 MMU.scala 126:29 MMU.scala 149:27]
  assign tlb_io_modify_pte_ppn_p2 = _T_81 ? 10'h0 : _GEN_86; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_ppn_p1 = _T_81 ? 10'h0 : _GEN_85; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_U = _T_81 ? 1'h0 : _GEN_80; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_X = _T_81 ? 1'h0 : _GEN_79; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_W = _T_81 ? 1'h0 : _GEN_78; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_R = _T_81 ? 1'h0 : _GEN_77; // @[MMU.scala 107:17 MMU.scala 150:27]
  assign tlb_io_modify_pte_V = _T_81 ? 1'h0 : _GEN_76; // @[MMU.scala 107:17 MMU.scala 150:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  csr_satp = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  csr_priv = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  csr_mxr = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  csr_sum = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  log_flush_one = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  log_flush_all = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  log_flush_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  status = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ptw_vpn_p2 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  ptw_vpn_p1 = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  _T_101 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _T_102 = _RAND_11[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      csr_satp <= 32'h0;
    end else if (ready) begin
      csr_satp <= io_csr_satp;
    end
    if (reset) begin
      csr_priv <= 2'h0;
    end else if (ready) begin
      csr_priv <= io_csr_priv;
    end
    if (reset) begin
      csr_mxr <= 1'h0;
    end else if (ready) begin
      csr_mxr <= io_csr_mxr;
    end
    if (reset) begin
      csr_sum <= 1'h0;
    end else if (ready) begin
      csr_sum <= io_csr_sum;
    end
    if (reset) begin
      log_flush_one <= 1'h0;
    end else if (_T_81) begin
      if (ready) begin
        log_flush_one <= 1'h0;
      end else if (_T_6) begin
        log_flush_one <= io_csr_flush_one;
      end
    end else if (_T_6) begin
      log_flush_one <= io_csr_flush_one;
    end
    if (reset) begin
      log_flush_all <= 1'h0;
    end else if (_T_81) begin
      if (ready) begin
        log_flush_all <= 1'h0;
      end else if (_T_6) begin
        log_flush_all <= io_csr_flush_all;
      end
    end else if (_T_6) begin
      log_flush_all <= io_csr_flush_all;
    end
    if (reset) begin
      log_flush_addr <= 32'h0;
    end else if (_T_81) begin
      if (ready) begin
        log_flush_addr <= 32'h0;
      end else if (_T_6) begin
        log_flush_addr <= io_csr_flush_addr;
      end
    end else if (_T_6) begin
      log_flush_addr <= io_csr_flush_addr;
    end
    if (reset) begin
      status <= 1'h0;
    end else if (_T_81) begin
      status <= _GEN_35;
    end else if (status) begin
      if (ptw_io_rsp_valid) begin
        status <= 1'h0;
      end
    end
    if (reset) begin
      ptw_vpn_p2 <= 10'h0;
    end else if (_T_81) begin
      if (_T_93) begin
        ptw_vpn_p2 <= tlb_io_query2_req_bits_p2;
      end else if (_T_87) begin
        ptw_vpn_p2 <= tlb_io_query_req_bits_p2;
      end
    end
    if (reset) begin
      ptw_vpn_p1 <= 10'h0;
    end else if (_T_81) begin
      if (_T_93) begin
        ptw_vpn_p1 <= tlb_io_query2_req_bits_p1;
      end else if (_T_87) begin
        ptw_vpn_p1 <= tlb_io_query_req_bits_p1;
      end
    end
    _T_101 <= ptw_io_mem_addr;
    _T_102 <= ptw_io_mem_mode;
  end
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [11:0] io_id_addr,
  output [31:0] io_id_rdata,
  output [1:0]  io_id_prv,
  input         io_mem_wrCSROp_valid,
  input  [11:0] io_mem_wrCSROp_addr,
  input  [31:0] io_mem_wrCSROp_data,
  input         io_mem_excep_valid,
  input  [31:0] io_mem_excep_code,
  input  [31:0] io_mem_excep_value,
  input  [31:0] io_mem_excep_pc,
  input         io_mem_excep_valid_inst,
  output        io_mem_inter_valid,
  output [31:0] io_mem_inter_bits,
  output [31:0] io_mmu_satp,
  output        io_mmu_flush_one,
  output        io_mmu_flush_all,
  output [31:0] io_mmu_flush_addr,
  output [1:0]  io_mmu_priv,
  output        io_mmu_mxr,
  output        io_mmu_sum,
  output        io_flush,
  output [31:0] io_csrNewPc
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] csr [0:1023]; // @[CSR.scala 76:16]
  wire [31:0] csr__T_45_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_45_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_86_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_86_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_87_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_87_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_mtvec_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mtvec_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_stvec_data; // @[CSR.scala 76:16]
  wire [9:0] csr_stvec_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_utvec_data; // @[CSR.scala 76:16]
  wire [9:0] csr_utvec_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_medeleg_data; // @[CSR.scala 76:16]
  wire [9:0] csr_medeleg_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_mideleg_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mideleg_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_sedeleg_data; // @[CSR.scala 76:16]
  wire [9:0] csr_sedeleg_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_sideleg_data; // @[CSR.scala 76:16]
  wire [9:0] csr_sideleg_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_mie_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mie_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_mip_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mip_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_250_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_250_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_251_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_251_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_384_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_384_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_mepc_r_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mepc_r_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_sepc_r_data; // @[CSR.scala 76:16]
  wire [9:0] csr_sepc_r_addr; // @[CSR.scala 76:16]
  wire [31:0] csr_uepc_r_data; // @[CSR.scala 76:16]
  wire [9:0] csr_uepc_r_addr; // @[CSR.scala 76:16]
  wire [31:0] csr__T_1_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_1_addr; // @[CSR.scala 76:16]
  wire  csr__T_1_mask; // @[CSR.scala 76:16]
  wire  csr__T_1_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_2_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_2_addr; // @[CSR.scala 76:16]
  wire  csr__T_2_mask; // @[CSR.scala 76:16]
  wire  csr__T_2_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_3_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_3_addr; // @[CSR.scala 76:16]
  wire  csr__T_3_mask; // @[CSR.scala 76:16]
  wire  csr__T_3_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_4_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_4_addr; // @[CSR.scala 76:16]
  wire  csr__T_4_mask; // @[CSR.scala 76:16]
  wire  csr__T_4_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_5_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_5_addr; // @[CSR.scala 76:16]
  wire  csr__T_5_mask; // @[CSR.scala 76:16]
  wire  csr__T_5_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_6_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_6_addr; // @[CSR.scala 76:16]
  wire  csr__T_6_mask; // @[CSR.scala 76:16]
  wire  csr__T_6_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_7_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_7_addr; // @[CSR.scala 76:16]
  wire  csr__T_7_mask; // @[CSR.scala 76:16]
  wire  csr__T_7_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_8_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_8_addr; // @[CSR.scala 76:16]
  wire  csr__T_8_mask; // @[CSR.scala 76:16]
  wire  csr__T_8_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_9_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_9_addr; // @[CSR.scala 76:16]
  wire  csr__T_9_mask; // @[CSR.scala 76:16]
  wire  csr__T_9_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_10_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_10_addr; // @[CSR.scala 76:16]
  wire  csr__T_10_mask; // @[CSR.scala 76:16]
  wire  csr__T_10_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_11_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_11_addr; // @[CSR.scala 76:16]
  wire  csr__T_11_mask; // @[CSR.scala 76:16]
  wire  csr__T_11_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_12_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_12_addr; // @[CSR.scala 76:16]
  wire  csr__T_12_mask; // @[CSR.scala 76:16]
  wire  csr__T_12_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_13_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_13_addr; // @[CSR.scala 76:16]
  wire  csr__T_13_mask; // @[CSR.scala 76:16]
  wire  csr__T_13_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_14_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_14_addr; // @[CSR.scala 76:16]
  wire  csr__T_14_mask; // @[CSR.scala 76:16]
  wire  csr__T_14_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_15_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_15_addr; // @[CSR.scala 76:16]
  wire  csr__T_15_mask; // @[CSR.scala 76:16]
  wire  csr__T_15_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_16_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_16_addr; // @[CSR.scala 76:16]
  wire  csr__T_16_mask; // @[CSR.scala 76:16]
  wire  csr__T_16_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_17_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_17_addr; // @[CSR.scala 76:16]
  wire  csr__T_17_mask; // @[CSR.scala 76:16]
  wire  csr__T_17_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_18_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_18_addr; // @[CSR.scala 76:16]
  wire  csr__T_18_mask; // @[CSR.scala 76:16]
  wire  csr__T_18_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_19_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_19_addr; // @[CSR.scala 76:16]
  wire  csr__T_19_mask; // @[CSR.scala 76:16]
  wire  csr__T_19_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_20_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_20_addr; // @[CSR.scala 76:16]
  wire  csr__T_20_mask; // @[CSR.scala 76:16]
  wire  csr__T_20_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_21_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_21_addr; // @[CSR.scala 76:16]
  wire  csr__T_21_mask; // @[CSR.scala 76:16]
  wire  csr__T_21_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_22_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_22_addr; // @[CSR.scala 76:16]
  wire  csr__T_22_mask; // @[CSR.scala 76:16]
  wire  csr__T_22_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_23_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_23_addr; // @[CSR.scala 76:16]
  wire  csr__T_23_mask; // @[CSR.scala 76:16]
  wire  csr__T_23_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_24_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_24_addr; // @[CSR.scala 76:16]
  wire  csr__T_24_mask; // @[CSR.scala 76:16]
  wire  csr__T_24_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_25_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_25_addr; // @[CSR.scala 76:16]
  wire  csr__T_25_mask; // @[CSR.scala 76:16]
  wire  csr__T_25_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_26_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_26_addr; // @[CSR.scala 76:16]
  wire  csr__T_26_mask; // @[CSR.scala 76:16]
  wire  csr__T_26_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_27_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_27_addr; // @[CSR.scala 76:16]
  wire  csr__T_27_mask; // @[CSR.scala 76:16]
  wire  csr__T_27_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_28_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_28_addr; // @[CSR.scala 76:16]
  wire  csr__T_28_mask; // @[CSR.scala 76:16]
  wire  csr__T_28_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_29_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_29_addr; // @[CSR.scala 76:16]
  wire  csr__T_29_mask; // @[CSR.scala 76:16]
  wire  csr__T_29_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_30_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_30_addr; // @[CSR.scala 76:16]
  wire  csr__T_30_mask; // @[CSR.scala 76:16]
  wire  csr__T_30_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_31_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_31_addr; // @[CSR.scala 76:16]
  wire  csr__T_31_mask; // @[CSR.scala 76:16]
  wire  csr__T_31_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_32_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_32_addr; // @[CSR.scala 76:16]
  wire  csr__T_32_mask; // @[CSR.scala 76:16]
  wire  csr__T_32_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_33_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_33_addr; // @[CSR.scala 76:16]
  wire  csr__T_33_mask; // @[CSR.scala 76:16]
  wire  csr__T_33_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_34_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_34_addr; // @[CSR.scala 76:16]
  wire  csr__T_34_mask; // @[CSR.scala 76:16]
  wire  csr__T_34_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_35_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_35_addr; // @[CSR.scala 76:16]
  wire  csr__T_35_mask; // @[CSR.scala 76:16]
  wire  csr__T_35_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_36_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_36_addr; // @[CSR.scala 76:16]
  wire  csr__T_36_mask; // @[CSR.scala 76:16]
  wire  csr__T_36_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_37_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_37_addr; // @[CSR.scala 76:16]
  wire  csr__T_37_mask; // @[CSR.scala 76:16]
  wire  csr__T_37_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_38_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_38_addr; // @[CSR.scala 76:16]
  wire  csr__T_38_mask; // @[CSR.scala 76:16]
  wire  csr__T_38_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_39_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_39_addr; // @[CSR.scala 76:16]
  wire  csr__T_39_mask; // @[CSR.scala 76:16]
  wire  csr__T_39_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_40_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_40_addr; // @[CSR.scala 76:16]
  wire  csr__T_40_mask; // @[CSR.scala 76:16]
  wire  csr__T_40_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_119_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_119_addr; // @[CSR.scala 76:16]
  wire  csr__T_119_mask; // @[CSR.scala 76:16]
  wire  csr__T_119_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_121_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_121_addr; // @[CSR.scala 76:16]
  wire  csr__T_121_mask; // @[CSR.scala 76:16]
  wire  csr__T_121_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_123_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_123_addr; // @[CSR.scala 76:16]
  wire  csr__T_123_mask; // @[CSR.scala 76:16]
  wire  csr__T_123_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_125_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_125_addr; // @[CSR.scala 76:16]
  wire  csr__T_125_mask; // @[CSR.scala 76:16]
  wire  csr__T_125_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_127_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_127_addr; // @[CSR.scala 76:16]
  wire  csr__T_127_mask; // @[CSR.scala 76:16]
  wire  csr__T_127_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_129_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_129_addr; // @[CSR.scala 76:16]
  wire  csr__T_129_mask; // @[CSR.scala 76:16]
  wire  csr__T_129_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_131_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_131_addr; // @[CSR.scala 76:16]
  wire  csr__T_131_mask; // @[CSR.scala 76:16]
  wire  csr__T_131_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_133_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_133_addr; // @[CSR.scala 76:16]
  wire  csr__T_133_mask; // @[CSR.scala 76:16]
  wire  csr__T_133_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_135_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_135_addr; // @[CSR.scala 76:16]
  wire  csr__T_135_mask; // @[CSR.scala 76:16]
  wire  csr__T_135_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_137_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_137_addr; // @[CSR.scala 76:16]
  wire  csr__T_137_mask; // @[CSR.scala 76:16]
  wire  csr__T_137_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_139_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_139_addr; // @[CSR.scala 76:16]
  wire  csr__T_139_mask; // @[CSR.scala 76:16]
  wire  csr__T_139_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_141_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_141_addr; // @[CSR.scala 76:16]
  wire  csr__T_141_mask; // @[CSR.scala 76:16]
  wire  csr__T_141_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_143_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_143_addr; // @[CSR.scala 76:16]
  wire  csr__T_143_mask; // @[CSR.scala 76:16]
  wire  csr__T_143_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_145_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_145_addr; // @[CSR.scala 76:16]
  wire  csr__T_145_mask; // @[CSR.scala 76:16]
  wire  csr__T_145_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_147_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_147_addr; // @[CSR.scala 76:16]
  wire  csr__T_147_mask; // @[CSR.scala 76:16]
  wire  csr__T_147_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_149_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_149_addr; // @[CSR.scala 76:16]
  wire  csr__T_149_mask; // @[CSR.scala 76:16]
  wire  csr__T_149_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_151_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_151_addr; // @[CSR.scala 76:16]
  wire  csr__T_151_mask; // @[CSR.scala 76:16]
  wire  csr__T_151_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_153_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_153_addr; // @[CSR.scala 76:16]
  wire  csr__T_153_mask; // @[CSR.scala 76:16]
  wire  csr__T_153_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_155_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_155_addr; // @[CSR.scala 76:16]
  wire  csr__T_155_mask; // @[CSR.scala 76:16]
  wire  csr__T_155_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_157_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_157_addr; // @[CSR.scala 76:16]
  wire  csr__T_157_mask; // @[CSR.scala 76:16]
  wire  csr__T_157_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_159_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_159_addr; // @[CSR.scala 76:16]
  wire  csr__T_159_mask; // @[CSR.scala 76:16]
  wire  csr__T_159_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_161_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_161_addr; // @[CSR.scala 76:16]
  wire  csr__T_161_mask; // @[CSR.scala 76:16]
  wire  csr__T_161_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_163_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_163_addr; // @[CSR.scala 76:16]
  wire  csr__T_163_mask; // @[CSR.scala 76:16]
  wire  csr__T_163_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_165_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_165_addr; // @[CSR.scala 76:16]
  wire  csr__T_165_mask; // @[CSR.scala 76:16]
  wire  csr__T_165_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_167_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_167_addr; // @[CSR.scala 76:16]
  wire  csr__T_167_mask; // @[CSR.scala 76:16]
  wire  csr__T_167_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_169_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_169_addr; // @[CSR.scala 76:16]
  wire  csr__T_169_mask; // @[CSR.scala 76:16]
  wire  csr__T_169_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_171_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_171_addr; // @[CSR.scala 76:16]
  wire  csr__T_171_mask; // @[CSR.scala 76:16]
  wire  csr__T_171_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_173_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_173_addr; // @[CSR.scala 76:16]
  wire  csr__T_173_mask; // @[CSR.scala 76:16]
  wire  csr__T_173_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_175_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_175_addr; // @[CSR.scala 76:16]
  wire  csr__T_175_mask; // @[CSR.scala 76:16]
  wire  csr__T_175_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_177_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_177_addr; // @[CSR.scala 76:16]
  wire  csr__T_177_mask; // @[CSR.scala 76:16]
  wire  csr__T_177_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_179_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_179_addr; // @[CSR.scala 76:16]
  wire  csr__T_179_mask; // @[CSR.scala 76:16]
  wire  csr__T_179_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_181_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_181_addr; // @[CSR.scala 76:16]
  wire  csr__T_181_mask; // @[CSR.scala 76:16]
  wire  csr__T_181_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_183_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_183_addr; // @[CSR.scala 76:16]
  wire  csr__T_183_mask; // @[CSR.scala 76:16]
  wire  csr__T_183_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_185_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_185_addr; // @[CSR.scala 76:16]
  wire  csr__T_185_mask; // @[CSR.scala 76:16]
  wire  csr__T_185_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_187_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_187_addr; // @[CSR.scala 76:16]
  wire  csr__T_187_mask; // @[CSR.scala 76:16]
  wire  csr__T_187_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_189_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_189_addr; // @[CSR.scala 76:16]
  wire  csr__T_189_mask; // @[CSR.scala 76:16]
  wire  csr__T_189_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_191_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_191_addr; // @[CSR.scala 76:16]
  wire  csr__T_191_mask; // @[CSR.scala 76:16]
  wire  csr__T_191_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_193_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_193_addr; // @[CSR.scala 76:16]
  wire  csr__T_193_mask; // @[CSR.scala 76:16]
  wire  csr__T_193_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_195_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_195_addr; // @[CSR.scala 76:16]
  wire  csr__T_195_mask; // @[CSR.scala 76:16]
  wire  csr__T_195_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_197_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_197_addr; // @[CSR.scala 76:16]
  wire  csr__T_197_mask; // @[CSR.scala 76:16]
  wire  csr__T_197_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_247_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_247_addr; // @[CSR.scala 76:16]
  wire  csr__T_247_mask; // @[CSR.scala 76:16]
  wire  csr__T_247_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_249_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_249_addr; // @[CSR.scala 76:16]
  wire  csr__T_249_mask; // @[CSR.scala 76:16]
  wire  csr__T_249_en; // @[CSR.scala 76:16]
  wire [31:0] csr_mcause_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mcause_addr; // @[CSR.scala 76:16]
  wire  csr_mcause_mask; // @[CSR.scala 76:16]
  wire  csr_mcause_en; // @[CSR.scala 76:16]
  wire [31:0] csr_scause_data; // @[CSR.scala 76:16]
  wire [9:0] csr_scause_addr; // @[CSR.scala 76:16]
  wire  csr_scause_mask; // @[CSR.scala 76:16]
  wire  csr_scause_en; // @[CSR.scala 76:16]
  wire [31:0] csr_ucause_data; // @[CSR.scala 76:16]
  wire [9:0] csr_ucause_addr; // @[CSR.scala 76:16]
  wire  csr_ucause_mask; // @[CSR.scala 76:16]
  wire  csr_ucause_en; // @[CSR.scala 76:16]
  wire [31:0] csr_mtval_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mtval_addr; // @[CSR.scala 76:16]
  wire  csr_mtval_mask; // @[CSR.scala 76:16]
  wire  csr_mtval_en; // @[CSR.scala 76:16]
  wire [31:0] csr_stval_data; // @[CSR.scala 76:16]
  wire [9:0] csr_stval_addr; // @[CSR.scala 76:16]
  wire  csr_stval_mask; // @[CSR.scala 76:16]
  wire  csr_stval_en; // @[CSR.scala 76:16]
  wire [31:0] csr_utval_data; // @[CSR.scala 76:16]
  wire [9:0] csr_utval_addr; // @[CSR.scala 76:16]
  wire  csr_utval_mask; // @[CSR.scala 76:16]
  wire  csr_utval_en; // @[CSR.scala 76:16]
  wire [31:0] csr__T_257_data; // @[CSR.scala 76:16]
  wire [9:0] csr__T_257_addr; // @[CSR.scala 76:16]
  wire  csr__T_257_mask; // @[CSR.scala 76:16]
  wire  csr__T_257_en; // @[CSR.scala 76:16]
  wire [31:0] csr_mepc_w_data; // @[CSR.scala 76:16]
  wire [9:0] csr_mepc_w_addr; // @[CSR.scala 76:16]
  wire  csr_mepc_w_mask; // @[CSR.scala 76:16]
  wire  csr_mepc_w_en; // @[CSR.scala 76:16]
  wire [31:0] csr_sepc_w_data; // @[CSR.scala 76:16]
  wire [9:0] csr_sepc_w_addr; // @[CSR.scala 76:16]
  wire  csr_sepc_w_mask; // @[CSR.scala 76:16]
  wire  csr_sepc_w_en; // @[CSR.scala 76:16]
  wire [31:0] csr_uepc_w_data; // @[CSR.scala 76:16]
  wire [9:0] csr_uepc_w_addr; // @[CSR.scala 76:16]
  wire  csr_uepc_w_mask; // @[CSR.scala 76:16]
  wire  csr_uepc_w_en; // @[CSR.scala 76:16]
  reg [1:0] prv; // @[CSR.scala 20:24]
  reg  mstatus_SD; // @[CSR.scala 116:24]
  reg [7:0] mstatus_zero1; // @[CSR.scala 116:24]
  reg  mstatus_TSR; // @[CSR.scala 116:24]
  reg  mstatus_TW; // @[CSR.scala 116:24]
  reg  mstatus_TVM; // @[CSR.scala 116:24]
  reg  mstatus_MXR; // @[CSR.scala 116:24]
  reg  mstatus_SUM; // @[CSR.scala 116:24]
  reg  mstatus_MPriv; // @[CSR.scala 116:24]
  reg [1:0] mstatus_XS; // @[CSR.scala 116:24]
  reg [1:0] mstatus_FS; // @[CSR.scala 116:24]
  reg [1:0] mstatus_MPP; // @[CSR.scala 116:24]
  reg [1:0] mstatus_old_HPP; // @[CSR.scala 116:24]
  reg  mstatus_SPP; // @[CSR.scala 116:24]
  reg  mstatus_MPIE; // @[CSR.scala 116:24]
  reg  mstatus_old_HPIE; // @[CSR.scala 116:24]
  reg  mstatus_SPIE; // @[CSR.scala 116:24]
  reg  mstatus_UPIE; // @[CSR.scala 116:24]
  reg  mstatus_MIE; // @[CSR.scala 116:24]
  reg  mstatus_old_HIE; // @[CSR.scala 116:24]
  reg  mstatus_SIE; // @[CSR.scala 116:24]
  reg  mstatus_UIE; // @[CSR.scala 116:24]
  reg [63:0] mtime; // @[CSR.scala 117:22]
  wire [63:0] _T_43 = mtime + 64'h1; // @[CSR.scala 118:18]
  wire [10:0] _T_54 = {mstatus_old_HPP,mstatus_SPP,mstatus_MPIE,mstatus_old_HPIE,mstatus_SPIE,mstatus_UPIE,mstatus_MIE,mstatus_old_HIE,mstatus_SIE,mstatus_UIE}; // @[CSR.scala 131:29]
  wire [7:0] _T_58 = {mstatus_SUM,mstatus_MPriv,mstatus_XS,mstatus_FS,mstatus_MPP}; // @[CSR.scala 131:29]
  wire [31:0] _T_65 = {mstatus_SD,mstatus_zero1,mstatus_TSR,mstatus_TW,mstatus_TVM,mstatus_MXR,_T_58,_T_54}; // @[CSR.scala 131:29]
  wire  _T_92 = 12'hf11 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_93 = _T_92 ? 32'h91d : csr__T_45_data; // @[Mux.scala 80:57]
  wire  _T_94 = 12'hf12 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_95 = _T_94 ? 32'h8fffffff : _T_93; // @[Mux.scala 80:57]
  wire  _T_96 = 12'hf13 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_97 = _T_96 ? 32'h91d : _T_95; // @[Mux.scala 80:57]
  wire  _T_98 = 12'hf14 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_99 = _T_98 ? 32'h0 : _T_97; // @[Mux.scala 80:57]
  wire  _T_100 = 12'h301 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_101 = _T_100 ? 32'h40141100 : _T_99; // @[Mux.scala 80:57]
  wire  _T_102 = 12'h300 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_103 = _T_102 ? _T_65 : _T_101; // @[Mux.scala 80:57]
  wire  _T_104 = 12'h100 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_105 = _T_104 ? _T_65 : _T_103; // @[Mux.scala 80:57]
  wire  _T_106 = 12'h104 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_107 = _T_106 ? csr__T_86_data : _T_105; // @[Mux.scala 80:57]
  wire  _T_108 = 12'h144 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_109 = _T_108 ? csr__T_87_data : _T_107; // @[Mux.scala 80:57]
  wire  _T_110 = 12'hc01 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_111 = _T_110 ? mtime[31:0] : _T_109; // @[Mux.scala 80:57]
  wire  _T_112 = 12'hc81 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_113 = _T_112 ? mtime[63:32] : _T_111; // @[Mux.scala 80:57]
  wire  _T_114 = 12'hc00 == io_id_addr; // @[Mux.scala 80:60]
  wire [31:0] _T_115 = _T_114 ? mtime[31:0] : _T_113; // @[Mux.scala 80:57]
  wire  _T_116 = 12'hc80 == io_id_addr; // @[Mux.scala 80:60]
  wire  _T_118 = 12'hf11 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_120 = 12'hf12 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_122 = 12'hf13 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_124 = 12'hf14 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_126 = 12'h300 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_128 = 12'h301 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_130 = 12'h302 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_132 = 12'h303 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_134 = 12'h304 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_136 = 12'h305 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_138 = 12'h306 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_140 = 12'h340 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_142 = 12'h341 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_144 = 12'h342 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_146 = 12'h343 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_148 = 12'h344 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_150 = 12'h100 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_152 = 12'h102 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_154 = 12'h103 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_156 = 12'h104 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_158 = 12'h105 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_160 = 12'h106 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_162 = 12'h140 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_164 = 12'h141 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_166 = 12'h142 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_168 = 12'h143 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_170 = 12'h144 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_172 = 12'h180 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_174 = 12'h5 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_176 = 12'h40 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_178 = 12'h41 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_180 = 12'h42 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_182 = 12'h43 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_184 = 12'h44 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_186 = 12'h321 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_188 = 12'h322 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_190 = 12'hc01 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_192 = 12'hc81 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_194 = 12'hc00 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_196 = 12'hc80 == io_mem_wrCSROp_addr; // @[CSR.scala 145:14]
  wire  _T_198 = io_mem_wrCSROp_addr == 12'h300; // @[CSR.scala 149:30]
  wire  _GEN_244 = _T_198 ? io_mem_wrCSROp_data[0] : mstatus_UIE; // @[CSR.scala 149:48]
  wire  _GEN_245 = _T_198 ? io_mem_wrCSROp_data[1] : mstatus_SIE; // @[CSR.scala 149:48]
  wire  _GEN_248 = _T_198 ? io_mem_wrCSROp_data[4] : mstatus_UPIE; // @[CSR.scala 149:48]
  wire  _GEN_249 = _T_198 ? io_mem_wrCSROp_data[5] : mstatus_SPIE; // @[CSR.scala 149:48]
  wire  _GEN_251 = _T_198 ? io_mem_wrCSROp_data[7] : mstatus_MPIE; // @[CSR.scala 149:48]
  wire  _GEN_252 = _T_198 ? io_mem_wrCSROp_data[8] : mstatus_SPP; // @[CSR.scala 149:48]
  wire  _T_222 = io_mem_wrCSROp_addr == 12'h100; // @[CSR.scala 152:30]
  wire  _GEN_265 = _T_222 ? io_mem_wrCSROp_data[0] : _GEN_244; // @[CSR.scala 152:48]
  wire  _GEN_266 = _T_222 ? io_mem_wrCSROp_data[1] : _GEN_245; // @[CSR.scala 152:48]
  wire  _GEN_269 = _T_222 ? io_mem_wrCSROp_data[4] : _GEN_248; // @[CSR.scala 152:48]
  wire  _GEN_270 = _T_222 ? io_mem_wrCSROp_data[5] : _GEN_249; // @[CSR.scala 152:48]
  wire  _GEN_272 = _T_222 ? io_mem_wrCSROp_data[7] : _GEN_251; // @[CSR.scala 152:48]
  wire  _GEN_273 = _T_222 ? io_mem_wrCSROp_data[8] : _GEN_252; // @[CSR.scala 152:48]
  wire  _T_246 = io_mem_wrCSROp_addr == 12'h104; // @[CSR.scala 155:30]
  wire  _T_248 = io_mem_wrCSROp_addr == 12'h144; // @[CSR.scala 158:30]
  wire  _GEN_496 = io_mem_wrCSROp_valid ? _GEN_265 : mstatus_UIE; // @[CSR.scala 143:30]
  wire  _GEN_497 = io_mem_wrCSROp_valid ? _GEN_266 : mstatus_SIE; // @[CSR.scala 143:30]
  wire  _GEN_500 = io_mem_wrCSROp_valid ? _GEN_269 : mstatus_UPIE; // @[CSR.scala 143:30]
  wire  _GEN_501 = io_mem_wrCSROp_valid ? _GEN_270 : mstatus_SPIE; // @[CSR.scala 143:30]
  wire  _GEN_503 = io_mem_wrCSROp_valid ? _GEN_272 : mstatus_MPIE; // @[CSR.scala 143:30]
  wire  _GEN_504 = io_mem_wrCSROp_valid ? _GEN_273 : mstatus_SPP; // @[CSR.scala 143:30]
  wire [63:0] mtimecmp = {csr__T_250_data,csr__T_251_data}; // @[Cat.scala 29:58]
  wire  _T_252 = 2'h3 == prv; // @[Mux.scala 80:60]
  wire  _T_253 = _T_252 & mstatus_MIE; // @[Mux.scala 80:57]
  wire  _T_254 = 2'h1 == prv; // @[Mux.scala 80:60]
  wire  _T_255 = _T_254 ? mstatus_SIE : _T_253; // @[Mux.scala 80:57]
  wire  _T_256 = 2'h0 == prv; // @[Mux.scala 80:60]
  wire  ie = _T_256 ? mstatus_UIE : _T_255; // @[Mux.scala 80:57]
  wire  time_inter = mtime >= mtimecmp; // @[CSR.scala 194:27]
  wire  _T_258 = prv == 2'h3; // @[CSR.scala 206:10]
  wire  _T_260 = prv == 2'h1; // @[CSR.scala 208:10]
  wire  _T_262 = prv == 2'h0; // @[CSR.scala 209:10]
  wire  _T_265 = _T_258 & time_inter; // @[CSR.scala 211:22]
  wire  _T_267 = _T_260 & time_inter; // @[CSR.scala 213:22]
  wire  _T_269 = _T_262 & time_inter; // @[CSR.scala 214:22]
  wire [7:0] _T_274 = {_T_265,1'h0,_T_267,_T_269,csr_mip_data[3:0]}; // @[Cat.scala 29:58]
  wire [31:0] ipie = csr_mip_data & csr_mie_data; // @[CSR.scala 218:18]
  wire [31:0] _T_280 = ~csr_mideleg_data; // @[CSR.scala 219:23]
  wire [31:0] ipie_m = ipie & _T_280; // @[CSR.scala 219:21]
  wire [31:0] ipie_s = ipie & csr_mideleg_data; // @[CSR.scala 220:21]
  wire [1:0] _T_301 = ipie_s[3] ? 2'h3 : {{1'd0}, ipie_s[1]}; // @[Mux.scala 47:69]
  wire [2:0] _T_302 = ipie_s[4] ? 3'h4 : {{1'd0}, _T_301}; // @[Mux.scala 47:69]
  wire [2:0] _T_303 = ipie_s[5] ? 3'h5 : _T_302; // @[Mux.scala 47:69]
  wire [2:0] _T_304 = ipie_s[7] ? 3'h7 : _T_303; // @[Mux.scala 47:69]
  wire [3:0] _T_305 = ipie_s[8] ? 4'h8 : {{1'd0}, _T_304}; // @[Mux.scala 47:69]
  wire [3:0] _T_306 = ipie_s[9] ? 4'h9 : _T_305; // @[Mux.scala 47:69]
  wire [3:0] _T_307 = ipie_s[11] ? 4'hb : _T_306; // @[Mux.scala 47:69]
  wire [3:0] _T_308 = ipie_m[0] ? 4'h0 : _T_307; // @[Mux.scala 47:69]
  wire [3:0] _T_309 = ipie_m[1] ? 4'h1 : _T_308; // @[Mux.scala 47:69]
  wire [3:0] _T_310 = ipie_m[3] ? 4'h3 : _T_309; // @[Mux.scala 47:69]
  wire [3:0] _T_311 = ipie_m[4] ? 4'h4 : _T_310; // @[Mux.scala 47:69]
  wire [3:0] _T_312 = ipie_m[5] ? 4'h5 : _T_311; // @[Mux.scala 47:69]
  wire [3:0] _T_313 = ipie_m[7] ? 4'h7 : _T_312; // @[Mux.scala 47:69]
  wire [3:0] _T_314 = ipie_m[8] ? 4'h8 : _T_313; // @[Mux.scala 47:69]
  wire [3:0] _T_315 = ipie_m[9] ? 4'h9 : _T_314; // @[Mux.scala 47:69]
  wire [3:0] ic = ipie_m[11] ? 4'hb : _T_315; // @[Mux.scala 47:69]
  wire [31:0] _T_316 = csr_mideleg_data >> ic; // @[CSR.scala 250:36]
  wire [1:0] inter_new_mode = _T_316[0] ? 2'h1 : 2'h3; // @[CSR.scala 250:27]
  wire  _T_318 = inter_new_mode > prv; // @[CSR.scala 251:38]
  wire  _T_319 = inter_new_mode == prv; // @[CSR.scala 251:65]
  wire  _T_320 = _T_319 & ie; // @[CSR.scala 251:74]
  wire  inter_enable = _T_318 | _T_320; // @[CSR.scala 251:45]
  wire  _T_321 = |ipie; // @[CSR.scala 257:46]
  wire [31:0] _GEN_653 = {{28'd0}, ic}; // @[CSR.scala 258:48]
  wire  have_excep = io_mem_excep_valid & io_mem_excep_valid_inst; // @[CSR.scala 261:39]
  wire  _T_326 = io_mem_excep_code[31:2] == 30'h4; // @[Const.scala 133:40]
  wire  _T_328 = 2'h3 == io_mem_excep_code[1:0]; // @[Conditional.scala 37:30]
  wire  _T_329 = 2'h1 == io_mem_excep_code[1:0]; // @[Conditional.scala 37:30]
  wire  _T_330 = 2'h0 == io_mem_excep_code[1:0]; // @[Conditional.scala 37:30]
  wire  _GEN_528 = _T_330 | _GEN_500; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_529 = _T_330 ? 2'h0 : prv; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_530 = _T_330 ? csr_uepc_r_data : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_532 = _T_329 | _GEN_501; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_534 = _T_329 ? {{1'd0}, mstatus_SPP} : _GEN_529; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_535 = _T_329 ? csr_sepc_r_data : _GEN_530; // @[Conditional.scala 39:67]
  wire  _GEN_539 = _T_328 | _GEN_503; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_541 = _T_328 ? mstatus_MPP : _GEN_534; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_542 = _T_328 ? csr_mepc_r_data : _GEN_535; // @[Conditional.scala 40:58]
  wire  _T_331 = io_mem_excep_code == 32'h14; // @[CSR.scala 297:29]
  wire  _T_332 = io_mem_excep_code == 32'h15; // @[CSR.scala 297:65]
  wire  _T_333 = _T_331 | _T_332; // @[CSR.scala 297:49]
  wire [31:0] _T_335 = io_mem_excep_pc + 32'h4; // @[CSR.scala 298:38]
  wire  _T_337 = ~io_mem_excep_code[31]; // @[CSR.scala 303:10]
  wire [31:0] _T_339 = csr_medeleg_data >> io_mem_excep_code[4:0]; // @[CSR.scala 303:32]
  wire  _T_341 = ~_T_339[0]; // @[CSR.scala 303:24]
  wire  _T_342 = _T_337 & _T_341; // @[CSR.scala 303:21]
  wire [31:0] _T_345 = csr_mideleg_data >> io_mem_excep_code[4:0]; // @[CSR.scala 304:32]
  wire  _T_347 = ~_T_345[0]; // @[CSR.scala 304:24]
  wire  _T_348 = io_mem_excep_code[31] & _T_347; // @[CSR.scala 304:21]
  wire [31:0] _T_352 = csr_sedeleg_data >> io_mem_excep_code[4:0]; // @[CSR.scala 305:32]
  wire  _T_354 = ~_T_352[0]; // @[CSR.scala 305:24]
  wire  _T_355 = _T_337 & _T_354; // @[CSR.scala 305:21]
  wire [31:0] _T_358 = csr_sideleg_data >> io_mem_excep_code[4:0]; // @[CSR.scala 306:32]
  wire  _T_360 = ~_T_358[0]; // @[CSR.scala 306:24]
  wire  _T_361 = io_mem_excep_code[31] & _T_360; // @[CSR.scala 306:21]
  wire [1:0] _T_362 = _T_361 ? 2'h1 : 2'h0; // @[Mux.scala 47:69]
  wire [1:0] _T_363 = _T_355 ? 2'h1 : _T_362; // @[Mux.scala 47:69]
  wire [1:0] _T_364 = _T_348 ? 2'h3 : _T_363; // @[Mux.scala 47:69]
  wire [1:0] _T_365 = _T_342 ? 2'h3 : _T_364; // @[Mux.scala 47:69]
  wire [1:0] _GEN_588 = _T_333 ? prv : _T_365; // @[CSR.scala 297:86]
  wire [1:0] _GEN_612 = _T_326 ? _GEN_541 : _GEN_588; // @[CSR.scala 270:30]
  wire [1:0] nextPrv = have_excep ? _GEN_612 : prv; // @[CSR.scala 268:20]
  wire  _T_366 = 2'h3 == nextPrv; // @[Conditional.scala 37:30]
  wire  _T_367 = 2'h1 == nextPrv; // @[Conditional.scala 37:30]
  wire  _T_369 = 2'h0 == nextPrv; // @[Conditional.scala 37:30]
  wire  _GEN_564 = _T_367 ? 1'h0 : _T_369; // @[Conditional.scala 39:67]
  wire  _GEN_578 = _T_366 ? 1'h0 : _T_367; // @[Conditional.scala 40:58]
  wire  _GEN_584 = _T_366 ? 1'h0 : _GEN_564; // @[Conditional.scala 40:58]
  wire [31:0] _T_371 = _T_366 ? csr_mtvec_data : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _T_373 = _T_367 ? csr_stvec_data : _T_371; // @[Mux.scala 80:57]
  wire [31:0] _T_375 = _T_369 ? csr_utvec_data : _T_373; // @[Mux.scala 80:57]
  wire [31:0] _T_377 = {_T_375[31:2],2'h0}; // @[Cat.scala 29:58]
  wire  _T_379 = _T_375[1:0] == 2'h0; // @[CSR.scala 341:37]
  wire [34:0] _T_380 = 32'h4 * io_mem_excep_code; // @[CSR.scala 343:20]
  wire [34:0] _GEN_654 = {{3'd0}, _T_377}; // @[CSR.scala 343:14]
  wire [34:0] _T_382 = _GEN_654 + _T_380; // @[CSR.scala 343:14]
  wire [34:0] _T_383 = _T_379 ? {{3'd0}, _T_377} : _T_382; // @[CSR.scala 341:25]
  wire [34:0] _GEN_587 = _T_333 ? {{3'd0}, _T_335} : _T_383; // @[CSR.scala 297:86]
  wire  _GEN_593 = _T_333 ? 1'h0 : _T_366; // @[CSR.scala 297:86]
  wire  _GEN_600 = _T_333 ? 1'h0 : _GEN_578; // @[CSR.scala 297:86]
  wire  _GEN_606 = _T_333 ? 1'h0 : _GEN_584; // @[CSR.scala 297:86]
  wire [34:0] _GEN_613 = _T_326 ? {{3'd0}, _GEN_542} : _GEN_587; // @[CSR.scala 270:30]
  wire  _GEN_620 = _T_326 ? 1'h0 : _GEN_593; // @[CSR.scala 270:30]
  wire  _GEN_624 = _T_326 ? 1'h0 : _GEN_600; // @[CSR.scala 270:30]
  wire  _GEN_628 = _T_326 ? 1'h0 : _GEN_606; // @[CSR.scala 270:30]
  wire [34:0] _GEN_635 = have_excep ? _GEN_613 : 35'h0; // @[CSR.scala 268:20]
  wire  _GEN_642 = have_excep & _GEN_620; // @[CSR.scala 268:20]
  wire  _GEN_646 = have_excep & _GEN_624; // @[CSR.scala 268:20]
  wire  _GEN_650 = have_excep & _GEN_628; // @[CSR.scala 268:20]
  assign csr__T_45_addr = io_id_addr[9:0];
  assign csr__T_45_data = csr[csr__T_45_addr]; // @[CSR.scala 76:16]
  assign csr__T_86_addr = 10'h304;
  assign csr__T_86_data = csr[csr__T_86_addr]; // @[CSR.scala 76:16]
  assign csr__T_87_addr = 10'h344;
  assign csr__T_87_data = csr[csr__T_87_addr]; // @[CSR.scala 76:16]
  assign csr_mtvec_addr = 10'h305;
  assign csr_mtvec_data = csr[csr_mtvec_addr]; // @[CSR.scala 76:16]
  assign csr_stvec_addr = 10'h105;
  assign csr_stvec_data = csr[csr_stvec_addr]; // @[CSR.scala 76:16]
  assign csr_utvec_addr = 10'h5;
  assign csr_utvec_data = csr[csr_utvec_addr]; // @[CSR.scala 76:16]
  assign csr_medeleg_addr = 10'h302;
  assign csr_medeleg_data = csr[csr_medeleg_addr]; // @[CSR.scala 76:16]
  assign csr_mideleg_addr = 10'h303;
  assign csr_mideleg_data = csr[csr_mideleg_addr]; // @[CSR.scala 76:16]
  assign csr_sedeleg_addr = 10'h102;
  assign csr_sedeleg_data = csr[csr_sedeleg_addr]; // @[CSR.scala 76:16]
  assign csr_sideleg_addr = 10'h103;
  assign csr_sideleg_data = csr[csr_sideleg_addr]; // @[CSR.scala 76:16]
  assign csr_mie_addr = 10'h304;
  assign csr_mie_data = csr[csr_mie_addr]; // @[CSR.scala 76:16]
  assign csr_mip_addr = 10'h344;
  assign csr_mip_data = csr[csr_mip_addr]; // @[CSR.scala 76:16]
  assign csr__T_250_addr = 10'h322;
  assign csr__T_250_data = csr[csr__T_250_addr]; // @[CSR.scala 76:16]
  assign csr__T_251_addr = 10'h321;
  assign csr__T_251_data = csr[csr__T_251_addr]; // @[CSR.scala 76:16]
  assign csr__T_384_addr = 10'h180;
  assign csr__T_384_data = csr[csr__T_384_addr]; // @[CSR.scala 76:16]
  assign csr_mepc_r_addr = 10'h341;
  assign csr_mepc_r_data = csr[csr_mepc_r_addr]; // @[CSR.scala 76:16]
  assign csr_sepc_r_addr = 10'h141;
  assign csr_sepc_r_data = csr[csr_sepc_r_addr]; // @[CSR.scala 76:16]
  assign csr_uepc_r_addr = 10'h41;
  assign csr_uepc_r_data = csr[csr_uepc_r_addr]; // @[CSR.scala 76:16]
  assign csr__T_1_data = 32'h0;
  assign csr__T_1_addr = 10'h311;
  assign csr__T_1_mask = 1'h1;
  assign csr__T_1_en = reset;
  assign csr__T_2_data = 32'h0;
  assign csr__T_2_addr = 10'h312;
  assign csr__T_2_mask = 1'h1;
  assign csr__T_2_en = reset;
  assign csr__T_3_data = 32'h0;
  assign csr__T_3_addr = 10'h313;
  assign csr__T_3_mask = 1'h1;
  assign csr__T_3_en = reset;
  assign csr__T_4_data = 32'h0;
  assign csr__T_4_addr = 10'h314;
  assign csr__T_4_mask = 1'h1;
  assign csr__T_4_en = reset;
  assign csr__T_5_data = 32'h0;
  assign csr__T_5_addr = 10'h300;
  assign csr__T_5_mask = 1'h1;
  assign csr__T_5_en = reset;
  assign csr__T_6_data = 32'h0;
  assign csr__T_6_addr = 10'h301;
  assign csr__T_6_mask = 1'h1;
  assign csr__T_6_en = reset;
  assign csr__T_7_data = 32'h0;
  assign csr__T_7_addr = 10'h302;
  assign csr__T_7_mask = 1'h1;
  assign csr__T_7_en = reset;
  assign csr__T_8_data = 32'h0;
  assign csr__T_8_addr = 10'h303;
  assign csr__T_8_mask = 1'h1;
  assign csr__T_8_en = reset;
  assign csr__T_9_data = 32'h0;
  assign csr__T_9_addr = 10'h304;
  assign csr__T_9_mask = 1'h1;
  assign csr__T_9_en = reset;
  assign csr__T_10_data = 32'h0;
  assign csr__T_10_addr = 10'h305;
  assign csr__T_10_mask = 1'h1;
  assign csr__T_10_en = reset;
  assign csr__T_11_data = 32'h0;
  assign csr__T_11_addr = 10'h306;
  assign csr__T_11_mask = 1'h1;
  assign csr__T_11_en = reset;
  assign csr__T_12_data = 32'h0;
  assign csr__T_12_addr = 10'h340;
  assign csr__T_12_mask = 1'h1;
  assign csr__T_12_en = reset;
  assign csr__T_13_data = 32'h0;
  assign csr__T_13_addr = 10'h341;
  assign csr__T_13_mask = 1'h1;
  assign csr__T_13_en = reset;
  assign csr__T_14_data = 32'h0;
  assign csr__T_14_addr = 10'h342;
  assign csr__T_14_mask = 1'h1;
  assign csr__T_14_en = reset;
  assign csr__T_15_data = 32'h0;
  assign csr__T_15_addr = 10'h343;
  assign csr__T_15_mask = 1'h1;
  assign csr__T_15_en = reset;
  assign csr__T_16_data = 32'h0;
  assign csr__T_16_addr = 10'h344;
  assign csr__T_16_mask = 1'h1;
  assign csr__T_16_en = reset;
  assign csr__T_17_data = 32'h0;
  assign csr__T_17_addr = 10'h100;
  assign csr__T_17_mask = 1'h1;
  assign csr__T_17_en = reset;
  assign csr__T_18_data = 32'h0;
  assign csr__T_18_addr = 10'h102;
  assign csr__T_18_mask = 1'h1;
  assign csr__T_18_en = reset;
  assign csr__T_19_data = 32'h0;
  assign csr__T_19_addr = 10'h103;
  assign csr__T_19_mask = 1'h1;
  assign csr__T_19_en = reset;
  assign csr__T_20_data = 32'h0;
  assign csr__T_20_addr = 10'h104;
  assign csr__T_20_mask = 1'h1;
  assign csr__T_20_en = reset;
  assign csr__T_21_data = 32'h0;
  assign csr__T_21_addr = 10'h105;
  assign csr__T_21_mask = 1'h1;
  assign csr__T_21_en = reset;
  assign csr__T_22_data = 32'h0;
  assign csr__T_22_addr = 10'h106;
  assign csr__T_22_mask = 1'h1;
  assign csr__T_22_en = reset;
  assign csr__T_23_data = 32'h0;
  assign csr__T_23_addr = 10'h140;
  assign csr__T_23_mask = 1'h1;
  assign csr__T_23_en = reset;
  assign csr__T_24_data = 32'h0;
  assign csr__T_24_addr = 10'h141;
  assign csr__T_24_mask = 1'h1;
  assign csr__T_24_en = reset;
  assign csr__T_25_data = 32'h0;
  assign csr__T_25_addr = 10'h142;
  assign csr__T_25_mask = 1'h1;
  assign csr__T_25_en = reset;
  assign csr__T_26_data = 32'h0;
  assign csr__T_26_addr = 10'h143;
  assign csr__T_26_mask = 1'h1;
  assign csr__T_26_en = reset;
  assign csr__T_27_data = 32'h0;
  assign csr__T_27_addr = 10'h144;
  assign csr__T_27_mask = 1'h1;
  assign csr__T_27_en = reset;
  assign csr__T_28_data = 32'h0;
  assign csr__T_28_addr = 10'h180;
  assign csr__T_28_mask = 1'h1;
  assign csr__T_28_en = reset;
  assign csr__T_29_data = 32'h0;
  assign csr__T_29_addr = 10'h5;
  assign csr__T_29_mask = 1'h1;
  assign csr__T_29_en = reset;
  assign csr__T_30_data = 32'h0;
  assign csr__T_30_addr = 10'h40;
  assign csr__T_30_mask = 1'h1;
  assign csr__T_30_en = reset;
  assign csr__T_31_data = 32'h0;
  assign csr__T_31_addr = 10'h41;
  assign csr__T_31_mask = 1'h1;
  assign csr__T_31_en = reset;
  assign csr__T_32_data = 32'h0;
  assign csr__T_32_addr = 10'h42;
  assign csr__T_32_mask = 1'h1;
  assign csr__T_32_en = reset;
  assign csr__T_33_data = 32'h0;
  assign csr__T_33_addr = 10'h43;
  assign csr__T_33_mask = 1'h1;
  assign csr__T_33_en = reset;
  assign csr__T_34_data = 32'h0;
  assign csr__T_34_addr = 10'h44;
  assign csr__T_34_mask = 1'h1;
  assign csr__T_34_en = reset;
  assign csr__T_35_data = 32'h0;
  assign csr__T_35_addr = 10'h321;
  assign csr__T_35_mask = 1'h1;
  assign csr__T_35_en = reset;
  assign csr__T_36_data = 32'h0;
  assign csr__T_36_addr = 10'h322;
  assign csr__T_36_mask = 1'h1;
  assign csr__T_36_en = reset;
  assign csr__T_37_data = 32'h0;
  assign csr__T_37_addr = 10'h1;
  assign csr__T_37_mask = 1'h1;
  assign csr__T_37_en = reset;
  assign csr__T_38_data = 32'h0;
  assign csr__T_38_addr = 10'h81;
  assign csr__T_38_mask = 1'h1;
  assign csr__T_38_en = reset;
  assign csr__T_39_data = 32'h0;
  assign csr__T_39_addr = 10'h0;
  assign csr__T_39_mask = 1'h1;
  assign csr__T_39_en = reset;
  assign csr__T_40_data = 32'h0;
  assign csr__T_40_addr = 10'h80;
  assign csr__T_40_mask = 1'h1;
  assign csr__T_40_en = reset;
  assign csr__T_119_data = io_mem_wrCSROp_data;
  assign csr__T_119_addr = 10'h311;
  assign csr__T_119_mask = 1'h1;
  assign csr__T_119_en = io_mem_wrCSROp_valid & _T_118;
  assign csr__T_121_data = io_mem_wrCSROp_data;
  assign csr__T_121_addr = 10'h312;
  assign csr__T_121_mask = 1'h1;
  assign csr__T_121_en = io_mem_wrCSROp_valid & _T_120;
  assign csr__T_123_data = io_mem_wrCSROp_data;
  assign csr__T_123_addr = 10'h313;
  assign csr__T_123_mask = 1'h1;
  assign csr__T_123_en = io_mem_wrCSROp_valid & _T_122;
  assign csr__T_125_data = io_mem_wrCSROp_data;
  assign csr__T_125_addr = 10'h314;
  assign csr__T_125_mask = 1'h1;
  assign csr__T_125_en = io_mem_wrCSROp_valid & _T_124;
  assign csr__T_127_data = io_mem_wrCSROp_data;
  assign csr__T_127_addr = 10'h300;
  assign csr__T_127_mask = 1'h1;
  assign csr__T_127_en = io_mem_wrCSROp_valid & _T_126;
  assign csr__T_129_data = io_mem_wrCSROp_data;
  assign csr__T_129_addr = 10'h301;
  assign csr__T_129_mask = 1'h1;
  assign csr__T_129_en = io_mem_wrCSROp_valid & _T_128;
  assign csr__T_131_data = io_mem_wrCSROp_data;
  assign csr__T_131_addr = 10'h302;
  assign csr__T_131_mask = 1'h1;
  assign csr__T_131_en = io_mem_wrCSROp_valid & _T_130;
  assign csr__T_133_data = io_mem_wrCSROp_data;
  assign csr__T_133_addr = 10'h303;
  assign csr__T_133_mask = 1'h1;
  assign csr__T_133_en = io_mem_wrCSROp_valid & _T_132;
  assign csr__T_135_data = io_mem_wrCSROp_data;
  assign csr__T_135_addr = 10'h304;
  assign csr__T_135_mask = 1'h1;
  assign csr__T_135_en = io_mem_wrCSROp_valid & _T_134;
  assign csr__T_137_data = io_mem_wrCSROp_data;
  assign csr__T_137_addr = 10'h305;
  assign csr__T_137_mask = 1'h1;
  assign csr__T_137_en = io_mem_wrCSROp_valid & _T_136;
  assign csr__T_139_data = io_mem_wrCSROp_data;
  assign csr__T_139_addr = 10'h306;
  assign csr__T_139_mask = 1'h1;
  assign csr__T_139_en = io_mem_wrCSROp_valid & _T_138;
  assign csr__T_141_data = io_mem_wrCSROp_data;
  assign csr__T_141_addr = 10'h340;
  assign csr__T_141_mask = 1'h1;
  assign csr__T_141_en = io_mem_wrCSROp_valid & _T_140;
  assign csr__T_143_data = io_mem_wrCSROp_data;
  assign csr__T_143_addr = 10'h341;
  assign csr__T_143_mask = 1'h1;
  assign csr__T_143_en = io_mem_wrCSROp_valid & _T_142;
  assign csr__T_145_data = io_mem_wrCSROp_data;
  assign csr__T_145_addr = 10'h342;
  assign csr__T_145_mask = 1'h1;
  assign csr__T_145_en = io_mem_wrCSROp_valid & _T_144;
  assign csr__T_147_data = io_mem_wrCSROp_data;
  assign csr__T_147_addr = 10'h343;
  assign csr__T_147_mask = 1'h1;
  assign csr__T_147_en = io_mem_wrCSROp_valid & _T_146;
  assign csr__T_149_data = io_mem_wrCSROp_data;
  assign csr__T_149_addr = 10'h344;
  assign csr__T_149_mask = 1'h1;
  assign csr__T_149_en = io_mem_wrCSROp_valid & _T_148;
  assign csr__T_151_data = io_mem_wrCSROp_data;
  assign csr__T_151_addr = 10'h100;
  assign csr__T_151_mask = 1'h1;
  assign csr__T_151_en = io_mem_wrCSROp_valid & _T_150;
  assign csr__T_153_data = io_mem_wrCSROp_data;
  assign csr__T_153_addr = 10'h102;
  assign csr__T_153_mask = 1'h1;
  assign csr__T_153_en = io_mem_wrCSROp_valid & _T_152;
  assign csr__T_155_data = io_mem_wrCSROp_data;
  assign csr__T_155_addr = 10'h103;
  assign csr__T_155_mask = 1'h1;
  assign csr__T_155_en = io_mem_wrCSROp_valid & _T_154;
  assign csr__T_157_data = io_mem_wrCSROp_data;
  assign csr__T_157_addr = 10'h104;
  assign csr__T_157_mask = 1'h1;
  assign csr__T_157_en = io_mem_wrCSROp_valid & _T_156;
  assign csr__T_159_data = io_mem_wrCSROp_data;
  assign csr__T_159_addr = 10'h105;
  assign csr__T_159_mask = 1'h1;
  assign csr__T_159_en = io_mem_wrCSROp_valid & _T_158;
  assign csr__T_161_data = io_mem_wrCSROp_data;
  assign csr__T_161_addr = 10'h106;
  assign csr__T_161_mask = 1'h1;
  assign csr__T_161_en = io_mem_wrCSROp_valid & _T_160;
  assign csr__T_163_data = io_mem_wrCSROp_data;
  assign csr__T_163_addr = 10'h140;
  assign csr__T_163_mask = 1'h1;
  assign csr__T_163_en = io_mem_wrCSROp_valid & _T_162;
  assign csr__T_165_data = io_mem_wrCSROp_data;
  assign csr__T_165_addr = 10'h141;
  assign csr__T_165_mask = 1'h1;
  assign csr__T_165_en = io_mem_wrCSROp_valid & _T_164;
  assign csr__T_167_data = io_mem_wrCSROp_data;
  assign csr__T_167_addr = 10'h142;
  assign csr__T_167_mask = 1'h1;
  assign csr__T_167_en = io_mem_wrCSROp_valid & _T_166;
  assign csr__T_169_data = io_mem_wrCSROp_data;
  assign csr__T_169_addr = 10'h143;
  assign csr__T_169_mask = 1'h1;
  assign csr__T_169_en = io_mem_wrCSROp_valid & _T_168;
  assign csr__T_171_data = io_mem_wrCSROp_data;
  assign csr__T_171_addr = 10'h144;
  assign csr__T_171_mask = 1'h1;
  assign csr__T_171_en = io_mem_wrCSROp_valid & _T_170;
  assign csr__T_173_data = io_mem_wrCSROp_data;
  assign csr__T_173_addr = 10'h180;
  assign csr__T_173_mask = 1'h1;
  assign csr__T_173_en = io_mem_wrCSROp_valid & _T_172;
  assign csr__T_175_data = io_mem_wrCSROp_data;
  assign csr__T_175_addr = 10'h5;
  assign csr__T_175_mask = 1'h1;
  assign csr__T_175_en = io_mem_wrCSROp_valid & _T_174;
  assign csr__T_177_data = io_mem_wrCSROp_data;
  assign csr__T_177_addr = 10'h40;
  assign csr__T_177_mask = 1'h1;
  assign csr__T_177_en = io_mem_wrCSROp_valid & _T_176;
  assign csr__T_179_data = io_mem_wrCSROp_data;
  assign csr__T_179_addr = 10'h41;
  assign csr__T_179_mask = 1'h1;
  assign csr__T_179_en = io_mem_wrCSROp_valid & _T_178;
  assign csr__T_181_data = io_mem_wrCSROp_data;
  assign csr__T_181_addr = 10'h42;
  assign csr__T_181_mask = 1'h1;
  assign csr__T_181_en = io_mem_wrCSROp_valid & _T_180;
  assign csr__T_183_data = io_mem_wrCSROp_data;
  assign csr__T_183_addr = 10'h43;
  assign csr__T_183_mask = 1'h1;
  assign csr__T_183_en = io_mem_wrCSROp_valid & _T_182;
  assign csr__T_185_data = io_mem_wrCSROp_data;
  assign csr__T_185_addr = 10'h44;
  assign csr__T_185_mask = 1'h1;
  assign csr__T_185_en = io_mem_wrCSROp_valid & _T_184;
  assign csr__T_187_data = io_mem_wrCSROp_data;
  assign csr__T_187_addr = 10'h321;
  assign csr__T_187_mask = 1'h1;
  assign csr__T_187_en = io_mem_wrCSROp_valid & _T_186;
  assign csr__T_189_data = io_mem_wrCSROp_data;
  assign csr__T_189_addr = 10'h322;
  assign csr__T_189_mask = 1'h1;
  assign csr__T_189_en = io_mem_wrCSROp_valid & _T_188;
  assign csr__T_191_data = io_mem_wrCSROp_data;
  assign csr__T_191_addr = 10'h1;
  assign csr__T_191_mask = 1'h1;
  assign csr__T_191_en = io_mem_wrCSROp_valid & _T_190;
  assign csr__T_193_data = io_mem_wrCSROp_data;
  assign csr__T_193_addr = 10'h81;
  assign csr__T_193_mask = 1'h1;
  assign csr__T_193_en = io_mem_wrCSROp_valid & _T_192;
  assign csr__T_195_data = io_mem_wrCSROp_data;
  assign csr__T_195_addr = 10'h0;
  assign csr__T_195_mask = 1'h1;
  assign csr__T_195_en = io_mem_wrCSROp_valid & _T_194;
  assign csr__T_197_data = io_mem_wrCSROp_data;
  assign csr__T_197_addr = 10'h80;
  assign csr__T_197_mask = 1'h1;
  assign csr__T_197_en = io_mem_wrCSROp_valid & _T_196;
  assign csr__T_247_data = io_mem_wrCSROp_data;
  assign csr__T_247_addr = 10'h304;
  assign csr__T_247_mask = 1'h1;
  assign csr__T_247_en = io_mem_wrCSROp_valid & _T_246;
  assign csr__T_249_data = io_mem_wrCSROp_data;
  assign csr__T_249_addr = 10'h344;
  assign csr__T_249_mask = 1'h1;
  assign csr__T_249_en = io_mem_wrCSROp_valid & _T_248;
  assign csr_mcause_data = io_mem_excep_code;
  assign csr_mcause_addr = 10'h342;
  assign csr_mcause_mask = have_excep & _GEN_620;
  assign csr_mcause_en = 1'h1;
  assign csr_scause_data = io_mem_excep_code;
  assign csr_scause_addr = 10'h142;
  assign csr_scause_mask = have_excep & _GEN_624;
  assign csr_scause_en = 1'h1;
  assign csr_ucause_data = io_mem_excep_code;
  assign csr_ucause_addr = 10'h42;
  assign csr_ucause_mask = have_excep & _GEN_628;
  assign csr_ucause_en = 1'h1;
  assign csr_mtval_data = io_mem_excep_value;
  assign csr_mtval_addr = 10'h343;
  assign csr_mtval_mask = have_excep & _GEN_620;
  assign csr_mtval_en = 1'h1;
  assign csr_stval_data = io_mem_excep_value;
  assign csr_stval_addr = 10'h143;
  assign csr_stval_mask = have_excep & _GEN_624;
  assign csr_stval_en = 1'h1;
  assign csr_utval_data = io_mem_excep_value;
  assign csr_utval_addr = 10'h43;
  assign csr_utval_mask = have_excep & _GEN_628;
  assign csr_utval_en = 1'h1;
  assign csr__T_257_data = {24'h0,_T_274};
  assign csr__T_257_addr = 10'h344;
  assign csr__T_257_mask = 1'h1;
  assign csr__T_257_en = 1'h1;
  assign csr_mepc_w_data = io_mem_excep_pc;
  assign csr_mepc_w_addr = 10'h341;
  assign csr_mepc_w_mask = have_excep & _GEN_620;
  assign csr_mepc_w_en = have_excep & _GEN_620;
  assign csr_sepc_w_data = io_mem_excep_pc;
  assign csr_sepc_w_addr = 10'h141;
  assign csr_sepc_w_mask = have_excep & _GEN_624;
  assign csr_sepc_w_en = have_excep & _GEN_624;
  assign csr_uepc_w_data = io_mem_excep_pc;
  assign csr_uepc_w_addr = 10'h41;
  assign csr_uepc_w_mask = have_excep & _GEN_628;
  assign csr_uepc_w_en = have_excep & _GEN_628;
  assign io_id_rdata = _T_116 ? mtime[63:32] : _T_115; // @[CSR.scala 125:15]
  assign io_id_prv = prv; // @[CSR.scala 140:13]
  assign io_mem_inter_valid = inter_enable & _T_321; // @[CSR.scala 257:22]
  assign io_mem_inter_bits = 32'h80000000 | _GEN_653; // @[CSR.scala 258:22]
  assign io_mmu_satp = csr__T_384_data; // @[CSR.scala 350:15]
  assign io_mmu_flush_one = io_mem_excep_valid & _T_331; // @[CSR.scala 353:20]
  assign io_mmu_flush_all = io_mem_excep_valid & _T_332; // @[CSR.scala 354:20]
  assign io_mmu_flush_addr = io_mem_excep_value; // @[CSR.scala 355:21]
  assign io_mmu_priv = have_excep ? _GEN_612 : prv; // @[CSR.scala 356:15]
  assign io_mmu_mxr = mstatus_MXR; // @[CSR.scala 352:14]
  assign io_mmu_sum = mstatus_SUM; // @[CSR.scala 351:14]
  assign io_flush = io_mem_excep_valid & io_mem_excep_valid_inst; // @[CSR.scala 264:12]
  assign io_csrNewPc = _GEN_635[31:0]; // @[CSR.scala 265:15 CSR.scala 281:23 CSR.scala 288:23 CSR.scala 294:23 CSR.scala 298:19 CSR.scala 341:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    csr[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  prv = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  mstatus_SD = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  mstatus_zero1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  mstatus_TSR = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mstatus_TW = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mstatus_TVM = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  mstatus_MXR = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mstatus_SUM = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mstatus_MPriv = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  mstatus_XS = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  mstatus_FS = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  mstatus_MPP = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  mstatus_old_HPP = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  mstatus_SPP = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  mstatus_MPIE = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  mstatus_old_HPIE = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  mstatus_SPIE = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  mstatus_UPIE = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  mstatus_MIE = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mstatus_old_HIE = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mstatus_SIE = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  mstatus_UIE = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  mtime = _RAND_23[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(csr__T_1_en & csr__T_1_mask) begin
      csr[csr__T_1_addr] <= csr__T_1_data; // @[CSR.scala 76:16]
    end
    if(csr__T_2_en & csr__T_2_mask) begin
      csr[csr__T_2_addr] <= csr__T_2_data; // @[CSR.scala 76:16]
    end
    if(csr__T_3_en & csr__T_3_mask) begin
      csr[csr__T_3_addr] <= csr__T_3_data; // @[CSR.scala 76:16]
    end
    if(csr__T_4_en & csr__T_4_mask) begin
      csr[csr__T_4_addr] <= csr__T_4_data; // @[CSR.scala 76:16]
    end
    if(csr__T_5_en & csr__T_5_mask) begin
      csr[csr__T_5_addr] <= csr__T_5_data; // @[CSR.scala 76:16]
    end
    if(csr__T_6_en & csr__T_6_mask) begin
      csr[csr__T_6_addr] <= csr__T_6_data; // @[CSR.scala 76:16]
    end
    if(csr__T_7_en & csr__T_7_mask) begin
      csr[csr__T_7_addr] <= csr__T_7_data; // @[CSR.scala 76:16]
    end
    if(csr__T_8_en & csr__T_8_mask) begin
      csr[csr__T_8_addr] <= csr__T_8_data; // @[CSR.scala 76:16]
    end
    if(csr__T_9_en & csr__T_9_mask) begin
      csr[csr__T_9_addr] <= csr__T_9_data; // @[CSR.scala 76:16]
    end
    if(csr__T_10_en & csr__T_10_mask) begin
      csr[csr__T_10_addr] <= csr__T_10_data; // @[CSR.scala 76:16]
    end
    if(csr__T_11_en & csr__T_11_mask) begin
      csr[csr__T_11_addr] <= csr__T_11_data; // @[CSR.scala 76:16]
    end
    if(csr__T_12_en & csr__T_12_mask) begin
      csr[csr__T_12_addr] <= csr__T_12_data; // @[CSR.scala 76:16]
    end
    if(csr__T_13_en & csr__T_13_mask) begin
      csr[csr__T_13_addr] <= csr__T_13_data; // @[CSR.scala 76:16]
    end
    if(csr__T_14_en & csr__T_14_mask) begin
      csr[csr__T_14_addr] <= csr__T_14_data; // @[CSR.scala 76:16]
    end
    if(csr__T_15_en & csr__T_15_mask) begin
      csr[csr__T_15_addr] <= csr__T_15_data; // @[CSR.scala 76:16]
    end
    if(csr__T_16_en & csr__T_16_mask) begin
      csr[csr__T_16_addr] <= csr__T_16_data; // @[CSR.scala 76:16]
    end
    if(csr__T_17_en & csr__T_17_mask) begin
      csr[csr__T_17_addr] <= csr__T_17_data; // @[CSR.scala 76:16]
    end
    if(csr__T_18_en & csr__T_18_mask) begin
      csr[csr__T_18_addr] <= csr__T_18_data; // @[CSR.scala 76:16]
    end
    if(csr__T_19_en & csr__T_19_mask) begin
      csr[csr__T_19_addr] <= csr__T_19_data; // @[CSR.scala 76:16]
    end
    if(csr__T_20_en & csr__T_20_mask) begin
      csr[csr__T_20_addr] <= csr__T_20_data; // @[CSR.scala 76:16]
    end
    if(csr__T_21_en & csr__T_21_mask) begin
      csr[csr__T_21_addr] <= csr__T_21_data; // @[CSR.scala 76:16]
    end
    if(csr__T_22_en & csr__T_22_mask) begin
      csr[csr__T_22_addr] <= csr__T_22_data; // @[CSR.scala 76:16]
    end
    if(csr__T_23_en & csr__T_23_mask) begin
      csr[csr__T_23_addr] <= csr__T_23_data; // @[CSR.scala 76:16]
    end
    if(csr__T_24_en & csr__T_24_mask) begin
      csr[csr__T_24_addr] <= csr__T_24_data; // @[CSR.scala 76:16]
    end
    if(csr__T_25_en & csr__T_25_mask) begin
      csr[csr__T_25_addr] <= csr__T_25_data; // @[CSR.scala 76:16]
    end
    if(csr__T_26_en & csr__T_26_mask) begin
      csr[csr__T_26_addr] <= csr__T_26_data; // @[CSR.scala 76:16]
    end
    if(csr__T_27_en & csr__T_27_mask) begin
      csr[csr__T_27_addr] <= csr__T_27_data; // @[CSR.scala 76:16]
    end
    if(csr__T_28_en & csr__T_28_mask) begin
      csr[csr__T_28_addr] <= csr__T_28_data; // @[CSR.scala 76:16]
    end
    if(csr__T_29_en & csr__T_29_mask) begin
      csr[csr__T_29_addr] <= csr__T_29_data; // @[CSR.scala 76:16]
    end
    if(csr__T_30_en & csr__T_30_mask) begin
      csr[csr__T_30_addr] <= csr__T_30_data; // @[CSR.scala 76:16]
    end
    if(csr__T_31_en & csr__T_31_mask) begin
      csr[csr__T_31_addr] <= csr__T_31_data; // @[CSR.scala 76:16]
    end
    if(csr__T_32_en & csr__T_32_mask) begin
      csr[csr__T_32_addr] <= csr__T_32_data; // @[CSR.scala 76:16]
    end
    if(csr__T_33_en & csr__T_33_mask) begin
      csr[csr__T_33_addr] <= csr__T_33_data; // @[CSR.scala 76:16]
    end
    if(csr__T_34_en & csr__T_34_mask) begin
      csr[csr__T_34_addr] <= csr__T_34_data; // @[CSR.scala 76:16]
    end
    if(csr__T_35_en & csr__T_35_mask) begin
      csr[csr__T_35_addr] <= csr__T_35_data; // @[CSR.scala 76:16]
    end
    if(csr__T_36_en & csr__T_36_mask) begin
      csr[csr__T_36_addr] <= csr__T_36_data; // @[CSR.scala 76:16]
    end
    if(csr__T_37_en & csr__T_37_mask) begin
      csr[csr__T_37_addr] <= csr__T_37_data; // @[CSR.scala 76:16]
    end
    if(csr__T_38_en & csr__T_38_mask) begin
      csr[csr__T_38_addr] <= csr__T_38_data; // @[CSR.scala 76:16]
    end
    if(csr__T_39_en & csr__T_39_mask) begin
      csr[csr__T_39_addr] <= csr__T_39_data; // @[CSR.scala 76:16]
    end
    if(csr__T_40_en & csr__T_40_mask) begin
      csr[csr__T_40_addr] <= csr__T_40_data; // @[CSR.scala 76:16]
    end
    if(csr__T_119_en & csr__T_119_mask) begin
      csr[csr__T_119_addr] <= csr__T_119_data; // @[CSR.scala 76:16]
    end
    if(csr__T_121_en & csr__T_121_mask) begin
      csr[csr__T_121_addr] <= csr__T_121_data; // @[CSR.scala 76:16]
    end
    if(csr__T_123_en & csr__T_123_mask) begin
      csr[csr__T_123_addr] <= csr__T_123_data; // @[CSR.scala 76:16]
    end
    if(csr__T_125_en & csr__T_125_mask) begin
      csr[csr__T_125_addr] <= csr__T_125_data; // @[CSR.scala 76:16]
    end
    if(csr__T_127_en & csr__T_127_mask) begin
      csr[csr__T_127_addr] <= csr__T_127_data; // @[CSR.scala 76:16]
    end
    if(csr__T_129_en & csr__T_129_mask) begin
      csr[csr__T_129_addr] <= csr__T_129_data; // @[CSR.scala 76:16]
    end
    if(csr__T_131_en & csr__T_131_mask) begin
      csr[csr__T_131_addr] <= csr__T_131_data; // @[CSR.scala 76:16]
    end
    if(csr__T_133_en & csr__T_133_mask) begin
      csr[csr__T_133_addr] <= csr__T_133_data; // @[CSR.scala 76:16]
    end
    if(csr__T_135_en & csr__T_135_mask) begin
      csr[csr__T_135_addr] <= csr__T_135_data; // @[CSR.scala 76:16]
    end
    if(csr__T_137_en & csr__T_137_mask) begin
      csr[csr__T_137_addr] <= csr__T_137_data; // @[CSR.scala 76:16]
    end
    if(csr__T_139_en & csr__T_139_mask) begin
      csr[csr__T_139_addr] <= csr__T_139_data; // @[CSR.scala 76:16]
    end
    if(csr__T_141_en & csr__T_141_mask) begin
      csr[csr__T_141_addr] <= csr__T_141_data; // @[CSR.scala 76:16]
    end
    if(csr__T_143_en & csr__T_143_mask) begin
      csr[csr__T_143_addr] <= csr__T_143_data; // @[CSR.scala 76:16]
    end
    if(csr__T_145_en & csr__T_145_mask) begin
      csr[csr__T_145_addr] <= csr__T_145_data; // @[CSR.scala 76:16]
    end
    if(csr__T_147_en & csr__T_147_mask) begin
      csr[csr__T_147_addr] <= csr__T_147_data; // @[CSR.scala 76:16]
    end
    if(csr__T_149_en & csr__T_149_mask) begin
      csr[csr__T_149_addr] <= csr__T_149_data; // @[CSR.scala 76:16]
    end
    if(csr__T_151_en & csr__T_151_mask) begin
      csr[csr__T_151_addr] <= csr__T_151_data; // @[CSR.scala 76:16]
    end
    if(csr__T_153_en & csr__T_153_mask) begin
      csr[csr__T_153_addr] <= csr__T_153_data; // @[CSR.scala 76:16]
    end
    if(csr__T_155_en & csr__T_155_mask) begin
      csr[csr__T_155_addr] <= csr__T_155_data; // @[CSR.scala 76:16]
    end
    if(csr__T_157_en & csr__T_157_mask) begin
      csr[csr__T_157_addr] <= csr__T_157_data; // @[CSR.scala 76:16]
    end
    if(csr__T_159_en & csr__T_159_mask) begin
      csr[csr__T_159_addr] <= csr__T_159_data; // @[CSR.scala 76:16]
    end
    if(csr__T_161_en & csr__T_161_mask) begin
      csr[csr__T_161_addr] <= csr__T_161_data; // @[CSR.scala 76:16]
    end
    if(csr__T_163_en & csr__T_163_mask) begin
      csr[csr__T_163_addr] <= csr__T_163_data; // @[CSR.scala 76:16]
    end
    if(csr__T_165_en & csr__T_165_mask) begin
      csr[csr__T_165_addr] <= csr__T_165_data; // @[CSR.scala 76:16]
    end
    if(csr__T_167_en & csr__T_167_mask) begin
      csr[csr__T_167_addr] <= csr__T_167_data; // @[CSR.scala 76:16]
    end
    if(csr__T_169_en & csr__T_169_mask) begin
      csr[csr__T_169_addr] <= csr__T_169_data; // @[CSR.scala 76:16]
    end
    if(csr__T_171_en & csr__T_171_mask) begin
      csr[csr__T_171_addr] <= csr__T_171_data; // @[CSR.scala 76:16]
    end
    if(csr__T_173_en & csr__T_173_mask) begin
      csr[csr__T_173_addr] <= csr__T_173_data; // @[CSR.scala 76:16]
    end
    if(csr__T_175_en & csr__T_175_mask) begin
      csr[csr__T_175_addr] <= csr__T_175_data; // @[CSR.scala 76:16]
    end
    if(csr__T_177_en & csr__T_177_mask) begin
      csr[csr__T_177_addr] <= csr__T_177_data; // @[CSR.scala 76:16]
    end
    if(csr__T_179_en & csr__T_179_mask) begin
      csr[csr__T_179_addr] <= csr__T_179_data; // @[CSR.scala 76:16]
    end
    if(csr__T_181_en & csr__T_181_mask) begin
      csr[csr__T_181_addr] <= csr__T_181_data; // @[CSR.scala 76:16]
    end
    if(csr__T_183_en & csr__T_183_mask) begin
      csr[csr__T_183_addr] <= csr__T_183_data; // @[CSR.scala 76:16]
    end
    if(csr__T_185_en & csr__T_185_mask) begin
      csr[csr__T_185_addr] <= csr__T_185_data; // @[CSR.scala 76:16]
    end
    if(csr__T_187_en & csr__T_187_mask) begin
      csr[csr__T_187_addr] <= csr__T_187_data; // @[CSR.scala 76:16]
    end
    if(csr__T_189_en & csr__T_189_mask) begin
      csr[csr__T_189_addr] <= csr__T_189_data; // @[CSR.scala 76:16]
    end
    if(csr__T_191_en & csr__T_191_mask) begin
      csr[csr__T_191_addr] <= csr__T_191_data; // @[CSR.scala 76:16]
    end
    if(csr__T_193_en & csr__T_193_mask) begin
      csr[csr__T_193_addr] <= csr__T_193_data; // @[CSR.scala 76:16]
    end
    if(csr__T_195_en & csr__T_195_mask) begin
      csr[csr__T_195_addr] <= csr__T_195_data; // @[CSR.scala 76:16]
    end
    if(csr__T_197_en & csr__T_197_mask) begin
      csr[csr__T_197_addr] <= csr__T_197_data; // @[CSR.scala 76:16]
    end
    if(csr__T_247_en & csr__T_247_mask) begin
      csr[csr__T_247_addr] <= csr__T_247_data; // @[CSR.scala 76:16]
    end
    if(csr__T_249_en & csr__T_249_mask) begin
      csr[csr__T_249_addr] <= csr__T_249_data; // @[CSR.scala 76:16]
    end
    if(csr_mcause_en & csr_mcause_mask) begin
      csr[csr_mcause_addr] <= csr_mcause_data; // @[CSR.scala 76:16]
    end
    if(csr_scause_en & csr_scause_mask) begin
      csr[csr_scause_addr] <= csr_scause_data; // @[CSR.scala 76:16]
    end
    if(csr_ucause_en & csr_ucause_mask) begin
      csr[csr_ucause_addr] <= csr_ucause_data; // @[CSR.scala 76:16]
    end
    if(csr_mtval_en & csr_mtval_mask) begin
      csr[csr_mtval_addr] <= csr_mtval_data; // @[CSR.scala 76:16]
    end
    if(csr_stval_en & csr_stval_mask) begin
      csr[csr_stval_addr] <= csr_stval_data; // @[CSR.scala 76:16]
    end
    if(csr_utval_en & csr_utval_mask) begin
      csr[csr_utval_addr] <= csr_utval_data; // @[CSR.scala 76:16]
    end
    if(csr__T_257_en & csr__T_257_mask) begin
      csr[csr__T_257_addr] <= csr__T_257_data; // @[CSR.scala 76:16]
    end
    if(csr_mepc_w_en & csr_mepc_w_mask) begin
      csr[csr_mepc_w_addr] <= csr_mepc_w_data; // @[CSR.scala 76:16]
    end
    if(csr_sepc_w_en & csr_sepc_w_mask) begin
      csr[csr_sepc_w_addr] <= csr_sepc_w_data; // @[CSR.scala 76:16]
    end
    if(csr_uepc_w_en & csr_uepc_w_mask) begin
      csr[csr_uepc_w_addr] <= csr_uepc_w_data; // @[CSR.scala 76:16]
    end
    if (reset) begin
      prv <= 2'h3;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          prv <= mstatus_MPP;
        end else if (_T_329) begin
          prv <= {{1'd0}, mstatus_SPP};
        end else if (_T_330) begin
          prv <= 2'h0;
        end
      end else if (!(_T_333)) begin
        if (_T_342) begin
          prv <= 2'h3;
        end else if (_T_348) begin
          prv <= 2'h3;
        end else if (_T_355) begin
          prv <= 2'h1;
        end else if (_T_361) begin
          prv <= 2'h1;
        end else begin
          prv <= 2'h0;
        end
      end
    end
    if (reset) begin
      mstatus_SD <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_SD <= io_mem_wrCSROp_data[31];
      end else if (_T_198) begin
        mstatus_SD <= io_mem_wrCSROp_data[31];
      end
    end
    if (reset) begin
      mstatus_zero1 <= 8'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_zero1 <= io_mem_wrCSROp_data[30:23];
      end else if (_T_198) begin
        mstatus_zero1 <= io_mem_wrCSROp_data[30:23];
      end
    end
    if (reset) begin
      mstatus_TSR <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_TSR <= io_mem_wrCSROp_data[22];
      end else if (_T_198) begin
        mstatus_TSR <= io_mem_wrCSROp_data[22];
      end
    end
    if (reset) begin
      mstatus_TW <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_TW <= io_mem_wrCSROp_data[21];
      end else if (_T_198) begin
        mstatus_TW <= io_mem_wrCSROp_data[21];
      end
    end
    if (reset) begin
      mstatus_TVM <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_TVM <= io_mem_wrCSROp_data[20];
      end else if (_T_198) begin
        mstatus_TVM <= io_mem_wrCSROp_data[20];
      end
    end
    if (reset) begin
      mstatus_MXR <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_MXR <= io_mem_wrCSROp_data[19];
      end else if (_T_198) begin
        mstatus_MXR <= io_mem_wrCSROp_data[19];
      end
    end
    if (reset) begin
      mstatus_SUM <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_SUM <= io_mem_wrCSROp_data[18];
      end else if (_T_198) begin
        mstatus_SUM <= io_mem_wrCSROp_data[18];
      end
    end
    if (reset) begin
      mstatus_MPriv <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_MPriv <= io_mem_wrCSROp_data[17];
      end else if (_T_198) begin
        mstatus_MPriv <= io_mem_wrCSROp_data[17];
      end
    end
    if (reset) begin
      mstatus_XS <= 2'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_XS <= io_mem_wrCSROp_data[16:15];
      end else if (_T_198) begin
        mstatus_XS <= io_mem_wrCSROp_data[16:15];
      end
    end
    if (reset) begin
      mstatus_FS <= 2'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_FS <= io_mem_wrCSROp_data[14:13];
      end else if (_T_198) begin
        mstatus_FS <= io_mem_wrCSROp_data[14:13];
      end
    end
    if (reset) begin
      mstatus_MPP <= 2'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          mstatus_MPP <= 2'h0;
        end else if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_MPP <= io_mem_wrCSROp_data[12:11];
          end else if (_T_198) begin
            mstatus_MPP <= io_mem_wrCSROp_data[12:11];
          end
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_MPP <= io_mem_wrCSROp_data[12:11];
          end else if (_T_198) begin
            mstatus_MPP <= io_mem_wrCSROp_data[12:11];
          end
        end
      end else if (_T_366) begin
        mstatus_MPP <= prv;
      end else if (io_mem_wrCSROp_valid) begin
        if (_T_222) begin
          mstatus_MPP <= io_mem_wrCSROp_data[12:11];
        end else if (_T_198) begin
          mstatus_MPP <= io_mem_wrCSROp_data[12:11];
        end
      end
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_MPP <= io_mem_wrCSROp_data[12:11];
      end else if (_T_198) begin
        mstatus_MPP <= io_mem_wrCSROp_data[12:11];
      end
    end
    if (reset) begin
      mstatus_old_HPP <= 2'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_old_HPP <= io_mem_wrCSROp_data[10:9];
      end else if (_T_198) begin
        mstatus_old_HPP <= io_mem_wrCSROp_data[10:9];
      end
    end
    if (reset) begin
      mstatus_SPP <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_SPP <= io_mem_wrCSROp_data[8];
            end else if (_T_198) begin
              mstatus_SPP <= io_mem_wrCSROp_data[8];
            end
          end
        end else if (_T_329) begin
          mstatus_SPP <= 1'h0;
        end else if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end else if (_T_198) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end else if (_T_198) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end
        end
      end else if (_T_366) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end else if (_T_198) begin
            mstatus_SPP <= io_mem_wrCSROp_data[8];
          end
        end
      end else if (_T_367) begin
        mstatus_SPP <= _T_260;
      end else begin
        mstatus_SPP <= _GEN_504;
      end
    end else begin
      mstatus_SPP <= _GEN_504;
    end
    if (reset) begin
      mstatus_MPIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        mstatus_MPIE <= _GEN_539;
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_MPIE <= io_mem_wrCSROp_data[7];
          end else if (_T_198) begin
            mstatus_MPIE <= io_mem_wrCSROp_data[7];
          end
        end
      end else if (_T_366) begin
        mstatus_MPIE <= mstatus_MIE;
      end else if (io_mem_wrCSROp_valid) begin
        if (_T_222) begin
          mstatus_MPIE <= io_mem_wrCSROp_data[7];
        end else if (_T_198) begin
          mstatus_MPIE <= io_mem_wrCSROp_data[7];
        end
      end
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_MPIE <= io_mem_wrCSROp_data[7];
      end else if (_T_198) begin
        mstatus_MPIE <= io_mem_wrCSROp_data[7];
      end
    end
    if (reset) begin
      mstatus_old_HPIE <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_old_HPIE <= io_mem_wrCSROp_data[6];
      end else if (_T_198) begin
        mstatus_old_HPIE <= io_mem_wrCSROp_data[6];
      end
    end
    if (reset) begin
      mstatus_SPIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_SPIE <= io_mem_wrCSROp_data[5];
            end else if (_T_198) begin
              mstatus_SPIE <= io_mem_wrCSROp_data[5];
            end
          end
        end else begin
          mstatus_SPIE <= _GEN_532;
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SPIE <= io_mem_wrCSROp_data[5];
          end else if (_T_198) begin
            mstatus_SPIE <= io_mem_wrCSROp_data[5];
          end
        end
      end else if (_T_366) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SPIE <= io_mem_wrCSROp_data[5];
          end else if (_T_198) begin
            mstatus_SPIE <= io_mem_wrCSROp_data[5];
          end
        end
      end else if (_T_367) begin
        mstatus_SPIE <= mstatus_SIE;
      end else if (io_mem_wrCSROp_valid) begin
        if (_T_222) begin
          mstatus_SPIE <= io_mem_wrCSROp_data[5];
        end else if (_T_198) begin
          mstatus_SPIE <= io_mem_wrCSROp_data[5];
        end
      end
    end else begin
      mstatus_SPIE <= _GEN_501;
    end
    if (reset) begin
      mstatus_UPIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_UPIE <= io_mem_wrCSROp_data[4];
            end else if (_T_198) begin
              mstatus_UPIE <= io_mem_wrCSROp_data[4];
            end
          end
        end else if (_T_329) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_UPIE <= io_mem_wrCSROp_data[4];
            end else if (_T_198) begin
              mstatus_UPIE <= io_mem_wrCSROp_data[4];
            end
          end
        end else begin
          mstatus_UPIE <= _GEN_528;
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_UPIE <= io_mem_wrCSROp_data[4];
          end else if (_T_198) begin
            mstatus_UPIE <= io_mem_wrCSROp_data[4];
          end
        end
      end else if (_T_366) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_UPIE <= io_mem_wrCSROp_data[4];
          end else if (_T_198) begin
            mstatus_UPIE <= io_mem_wrCSROp_data[4];
          end
        end
      end else if (_T_367) begin
        mstatus_UPIE <= _GEN_500;
      end else if (_T_369) begin
        mstatus_UPIE <= mstatus_UIE;
      end else begin
        mstatus_UPIE <= _GEN_500;
      end
    end else begin
      mstatus_UPIE <= _GEN_500;
    end
    if (reset) begin
      mstatus_MIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          mstatus_MIE <= mstatus_MPIE;
        end else if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_MIE <= io_mem_wrCSROp_data[3];
          end else if (_T_198) begin
            mstatus_MIE <= io_mem_wrCSROp_data[3];
          end
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_MIE <= io_mem_wrCSROp_data[3];
          end else if (_T_198) begin
            mstatus_MIE <= io_mem_wrCSROp_data[3];
          end
        end
      end else if (_T_366) begin
        mstatus_MIE <= 1'h0;
      end else if (io_mem_wrCSROp_valid) begin
        if (_T_222) begin
          mstatus_MIE <= io_mem_wrCSROp_data[3];
        end else if (_T_198) begin
          mstatus_MIE <= io_mem_wrCSROp_data[3];
        end
      end
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_MIE <= io_mem_wrCSROp_data[3];
      end else if (_T_198) begin
        mstatus_MIE <= io_mem_wrCSROp_data[3];
      end
    end
    if (reset) begin
      mstatus_old_HIE <= 1'h0;
    end else if (io_mem_wrCSROp_valid) begin
      if (_T_222) begin
        mstatus_old_HIE <= io_mem_wrCSROp_data[2];
      end else if (_T_198) begin
        mstatus_old_HIE <= io_mem_wrCSROp_data[2];
      end
    end
    if (reset) begin
      mstatus_SIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_SIE <= io_mem_wrCSROp_data[1];
            end else if (_T_198) begin
              mstatus_SIE <= io_mem_wrCSROp_data[1];
            end
          end
        end else if (_T_329) begin
          mstatus_SIE <= mstatus_SPIE;
        end else if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end else if (_T_198) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end else if (_T_198) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end
        end
      end else if (_T_366) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end else if (_T_198) begin
            mstatus_SIE <= io_mem_wrCSROp_data[1];
          end
        end
      end else if (_T_367) begin
        mstatus_SIE <= 1'h0;
      end else begin
        mstatus_SIE <= _GEN_497;
      end
    end else begin
      mstatus_SIE <= _GEN_497;
    end
    if (reset) begin
      mstatus_UIE <= 1'h0;
    end else if (have_excep) begin
      if (_T_326) begin
        if (_T_328) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_UIE <= io_mem_wrCSROp_data[0];
            end else if (_T_198) begin
              mstatus_UIE <= io_mem_wrCSROp_data[0];
            end
          end
        end else if (_T_329) begin
          if (io_mem_wrCSROp_valid) begin
            if (_T_222) begin
              mstatus_UIE <= io_mem_wrCSROp_data[0];
            end else if (_T_198) begin
              mstatus_UIE <= io_mem_wrCSROp_data[0];
            end
          end
        end else if (_T_330) begin
          mstatus_UIE <= mstatus_MPIE;
        end else if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_UIE <= io_mem_wrCSROp_data[0];
          end else if (_T_198) begin
            mstatus_UIE <= io_mem_wrCSROp_data[0];
          end
        end
      end else if (_T_333) begin
        if (io_mem_wrCSROp_valid) begin
          if (_T_222) begin
            mstatus_UIE <= io_mem_wrCSROp_data[0];
          end else if (_T_198) begin
            mstatus_UIE <= io_mem_wrCSROp_data[0];
          end
        end
      end else if (_T_366) begin
        mstatus_UIE <= _GEN_496;
      end else if (_T_367) begin
        mstatus_UIE <= _GEN_496;
      end else if (_T_369) begin
        mstatus_UIE <= 1'h0;
      end else begin
        mstatus_UIE <= _GEN_496;
      end
    end else begin
      mstatus_UIE <= _GEN_496;
    end
    if (reset) begin
      mtime <= 64'h0;
    end else begin
      mtime <= _T_43;
    end
  end
endmodule
module Core(
  input         clock,
  input         reset,
  output [31:0] io_dev_if__addr,
  output [3:0]  io_dev_if__mode,
  input  [31:0] io_dev_if__rdata,
  input         io_dev_if__ok,
  output [31:0] io_dev_mem_addr,
  output [3:0]  io_dev_mem_mode,
  output [31:0] io_dev_mem_wdata,
  input  [31:0] io_dev_mem_rdata,
  input         io_dev_mem_ok,
  output [31:0] io_debug_idex_aluOp_rd1,
  output [31:0] io_debug_idex_aluOp_rd2,
  output [4:0]  io_debug_idex_aluOp_opt,
  output [4:0]  io_debug_idex_wrRegOp_addr,
  output [31:0] io_debug_idex_wrRegOp_data,
  output        io_debug_idex_wrRegOp_rdy,
  output        io_debug_idex_wrCSROp_valid,
  output [11:0] io_debug_idex_wrCSROp_addr,
  output [31:0] io_debug_idex_wrCSROp_data,
  output [31:0] io_debug_idex_store_data,
  output        io_debug_idex_excep_valid,
  output [31:0] io_debug_idex_excep_code,
  output [31:0] io_debug_idex_excep_value,
  output [31:0] io_debug_idex_excep_pc,
  output        io_debug_idex_excep_valid_inst,
  output [31:0] io_debug_ifpc,
  output [31:0] io_debug_reg_0,
  output [31:0] io_debug_reg_1,
  output [31:0] io_debug_reg_2,
  output [31:0] io_debug_reg_3,
  output [31:0] io_debug_reg_4,
  output [31:0] io_debug_reg_5,
  output [31:0] io_debug_reg_6,
  output [31:0] io_debug_reg_7,
  output [31:0] io_debug_reg_8,
  output [31:0] io_debug_reg_9,
  output [31:0] io_debug_reg_10,
  output [31:0] io_debug_reg_11,
  output [31:0] io_debug_reg_12,
  output [31:0] io_debug_reg_13,
  output [31:0] io_debug_reg_14,
  output [31:0] io_debug_reg_15,
  output [31:0] io_debug_reg_16,
  output [31:0] io_debug_reg_17,
  output [31:0] io_debug_reg_18,
  output [31:0] io_debug_reg_19,
  output [31:0] io_debug_reg_20,
  output [31:0] io_debug_reg_21,
  output [31:0] io_debug_reg_22,
  output [31:0] io_debug_reg_23,
  output [31:0] io_debug_reg_24,
  output [31:0] io_debug_reg_25,
  output [31:0] io_debug_reg_26,
  output [31:0] io_debug_reg_27,
  output [31:0] io_debug_reg_28,
  output [31:0] io_debug_reg_29,
  output [31:0] io_debug_reg_30,
  output [31:0] io_debug_reg_31,
  output        io_debug_finish_pc_valid,
  output [31:0] io_debug_finish_pc_bits
);
  wire  iff__clock; // @[Core.scala 20:19]
  wire  iff__reset; // @[Core.scala 20:19]
  wire [31:0] iff__io_mmu_addr; // @[Core.scala 20:19]
  wire [3:0] iff__io_mmu_mode; // @[Core.scala 20:19]
  wire [31:0] iff__io_mmu_rdata; // @[Core.scala 20:19]
  wire  iff__io_mmu_ok; // @[Core.scala 20:19]
  wire  iff__io_mmu_pageFault; // @[Core.scala 20:19]
  wire [31:0] iff__io_id_inst; // @[Core.scala 20:19]
  wire  iff__io_id_excep_valid; // @[Core.scala 20:19]
  wire [31:0] iff__io_id_excep_code; // @[Core.scala 20:19]
  wire [31:0] iff__io_id_excep_value; // @[Core.scala 20:19]
  wire [31:0] iff__io_id_excep_pc; // @[Core.scala 20:19]
  wire  iff__io_id_excep_valid_inst; // @[Core.scala 20:19]
  wire  iff__io_id_branch_valid; // @[Core.scala 20:19]
  wire [31:0] iff__io_id_branch_bits; // @[Core.scala 20:19]
  wire  iff__io_id_ready; // @[Core.scala 20:19]
  wire  id_clock; // @[Core.scala 21:19]
  wire  id_reset; // @[Core.scala 21:19]
  wire [31:0] id_io_iff_inst; // @[Core.scala 21:19]
  wire  id_io_iff_excep_valid; // @[Core.scala 21:19]
  wire [31:0] id_io_iff_excep_code; // @[Core.scala 21:19]
  wire [31:0] id_io_iff_excep_value; // @[Core.scala 21:19]
  wire [31:0] id_io_iff_excep_pc; // @[Core.scala 21:19]
  wire  id_io_iff_excep_valid_inst; // @[Core.scala 21:19]
  wire  id_io_iff_branch_valid; // @[Core.scala 21:19]
  wire [31:0] id_io_iff_branch_bits; // @[Core.scala 21:19]
  wire  id_io_iff_ready; // @[Core.scala 21:19]
  wire [4:0] id_io_reg_read1_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_reg_read1_data; // @[Core.scala 21:19]
  wire [4:0] id_io_reg_read2_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_reg_read2_data; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_aluOp_rd1; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_aluOp_rd2; // @[Core.scala 21:19]
  wire [4:0] id_io_ex_aluOp_opt; // @[Core.scala 21:19]
  wire [4:0] id_io_ex_wrRegOp_addr; // @[Core.scala 21:19]
  wire  id_io_ex_wrCSROp_valid; // @[Core.scala 21:19]
  wire [11:0] id_io_ex_wrCSROp_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_wrCSROp_data; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_store_data; // @[Core.scala 21:19]
  wire  id_io_ex_excep_valid; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_excep_code; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_excep_value; // @[Core.scala 21:19]
  wire [31:0] id_io_ex_excep_pc; // @[Core.scala 21:19]
  wire  id_io_ex_excep_valid_inst; // @[Core.scala 21:19]
  wire  id_io_ex_ready; // @[Core.scala 21:19]
  wire [11:0] id_io_csr_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_csr_rdata; // @[Core.scala 21:19]
  wire [1:0] id_io_csr_prv; // @[Core.scala 21:19]
  wire  id_io_flush; // @[Core.scala 21:19]
  wire [4:0] id_io_exWrRegOp_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_exWrRegOp_data; // @[Core.scala 21:19]
  wire  id_io_exWrRegOp_rdy; // @[Core.scala 21:19]
  wire [4:0] id_io_memWrRegOp_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_memWrRegOp_data; // @[Core.scala 21:19]
  wire  id_io_exWrCSROp_valid; // @[Core.scala 21:19]
  wire [11:0] id_io_exWrCSROp_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_exWrCSROp_data; // @[Core.scala 21:19]
  wire  id_io_memWrCSROp_valid; // @[Core.scala 21:19]
  wire [11:0] id_io_memWrCSROp_addr; // @[Core.scala 21:19]
  wire [31:0] id_io_memWrCSROp_data; // @[Core.scala 21:19]
  wire  ex_clock; // @[Core.scala 22:19]
  wire  ex_reset; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_aluOp_rd1; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_aluOp_rd2; // @[Core.scala 22:19]
  wire [4:0] ex_io_id_aluOp_opt; // @[Core.scala 22:19]
  wire [4:0] ex_io_id_wrRegOp_addr; // @[Core.scala 22:19]
  wire  ex_io_id_wrCSROp_valid; // @[Core.scala 22:19]
  wire [11:0] ex_io_id_wrCSROp_addr; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_wrCSROp_data; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_store_data; // @[Core.scala 22:19]
  wire  ex_io_id_excep_valid; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_excep_code; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_excep_value; // @[Core.scala 22:19]
  wire [31:0] ex_io_id_excep_pc; // @[Core.scala 22:19]
  wire  ex_io_id_excep_valid_inst; // @[Core.scala 22:19]
  wire  ex_io_id_ready; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_ramOp_addr; // @[Core.scala 22:19]
  wire [3:0] ex_io_mem_ramOp_mode; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_ramOp_wdata; // @[Core.scala 22:19]
  wire [4:0] ex_io_mem_wrRegOp_addr; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_wrRegOp_data; // @[Core.scala 22:19]
  wire  ex_io_mem_wrRegOp_rdy; // @[Core.scala 22:19]
  wire  ex_io_mem_wrCSROp_valid; // @[Core.scala 22:19]
  wire [11:0] ex_io_mem_wrCSROp_addr; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_wrCSROp_data; // @[Core.scala 22:19]
  wire  ex_io_mem_excep_valid; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_excep_code; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_excep_value; // @[Core.scala 22:19]
  wire [31:0] ex_io_mem_excep_pc; // @[Core.scala 22:19]
  wire  ex_io_mem_excep_valid_inst; // @[Core.scala 22:19]
  wire  ex_io_mem_ready; // @[Core.scala 22:19]
  wire  ex_io_flush; // @[Core.scala 22:19]
  wire  mem_clock; // @[Core.scala 23:19]
  wire  mem_reset; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_ramOp_addr; // @[Core.scala 23:19]
  wire [3:0] mem_io_ex_ramOp_mode; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_ramOp_wdata; // @[Core.scala 23:19]
  wire [4:0] mem_io_ex_wrRegOp_addr; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_wrRegOp_data; // @[Core.scala 23:19]
  wire  mem_io_ex_wrCSROp_valid; // @[Core.scala 23:19]
  wire [11:0] mem_io_ex_wrCSROp_addr; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_wrCSROp_data; // @[Core.scala 23:19]
  wire  mem_io_ex_excep_valid; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_excep_code; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_excep_value; // @[Core.scala 23:19]
  wire [31:0] mem_io_ex_excep_pc; // @[Core.scala 23:19]
  wire  mem_io_ex_excep_valid_inst; // @[Core.scala 23:19]
  wire  mem_io_ex_ready; // @[Core.scala 23:19]
  wire [31:0] mem_io_mmu_addr; // @[Core.scala 23:19]
  wire [3:0] mem_io_mmu_mode; // @[Core.scala 23:19]
  wire [31:0] mem_io_mmu_wdata; // @[Core.scala 23:19]
  wire [31:0] mem_io_mmu_rdata; // @[Core.scala 23:19]
  wire  mem_io_mmu_ok; // @[Core.scala 23:19]
  wire  mem_io_mmu_pageFault; // @[Core.scala 23:19]
  wire  mem_io_csr_wrCSROp_valid; // @[Core.scala 23:19]
  wire [11:0] mem_io_csr_wrCSROp_addr; // @[Core.scala 23:19]
  wire [31:0] mem_io_csr_wrCSROp_data; // @[Core.scala 23:19]
  wire  mem_io_csr_excep_valid; // @[Core.scala 23:19]
  wire [31:0] mem_io_csr_excep_code; // @[Core.scala 23:19]
  wire [31:0] mem_io_csr_excep_value; // @[Core.scala 23:19]
  wire [31:0] mem_io_csr_excep_pc; // @[Core.scala 23:19]
  wire  mem_io_csr_excep_valid_inst; // @[Core.scala 23:19]
  wire  mem_io_csr_inter_valid; // @[Core.scala 23:19]
  wire [31:0] mem_io_csr_inter_bits; // @[Core.scala 23:19]
  wire [4:0] mem_io_reg_addr; // @[Core.scala 23:19]
  wire [31:0] mem_io_reg_data; // @[Core.scala 23:19]
  wire  mem_io_flush; // @[Core.scala 23:19]
  wire  reg__clock; // @[Core.scala 24:19]
  wire [4:0] reg__io_id_read1_addr; // @[Core.scala 24:19]
  wire [31:0] reg__io_id_read1_data; // @[Core.scala 24:19]
  wire [4:0] reg__io_id_read2_addr; // @[Core.scala 24:19]
  wire [31:0] reg__io_id_read2_data; // @[Core.scala 24:19]
  wire [4:0] reg__io_mem_addr; // @[Core.scala 24:19]
  wire [31:0] reg__io_mem_data; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_0; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_1; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_2; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_3; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_4; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_5; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_6; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_7; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_8; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_9; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_10; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_11; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_12; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_13; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_14; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_15; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_16; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_17; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_18; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_19; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_20; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_21; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_22; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_23; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_24; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_25; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_26; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_27; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_28; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_29; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_30; // @[Core.scala 24:19]
  wire [31:0] reg__io_log_31; // @[Core.scala 24:19]
  wire  mmu_clock; // @[Core.scala 25:19]
  wire  mmu_reset; // @[Core.scala 25:19]
  wire [31:0] mmu_io_iff_addr; // @[Core.scala 25:19]
  wire [3:0] mmu_io_iff_mode; // @[Core.scala 25:19]
  wire [31:0] mmu_io_iff_rdata; // @[Core.scala 25:19]
  wire  mmu_io_iff_ok; // @[Core.scala 25:19]
  wire  mmu_io_iff_pageFault; // @[Core.scala 25:19]
  wire [31:0] mmu_io_mem_addr; // @[Core.scala 25:19]
  wire [3:0] mmu_io_mem_mode; // @[Core.scala 25:19]
  wire [31:0] mmu_io_mem_wdata; // @[Core.scala 25:19]
  wire [31:0] mmu_io_mem_rdata; // @[Core.scala 25:19]
  wire  mmu_io_mem_ok; // @[Core.scala 25:19]
  wire  mmu_io_mem_pageFault; // @[Core.scala 25:19]
  wire [31:0] mmu_io_csr_satp; // @[Core.scala 25:19]
  wire  mmu_io_csr_flush_one; // @[Core.scala 25:19]
  wire  mmu_io_csr_flush_all; // @[Core.scala 25:19]
  wire [31:0] mmu_io_csr_flush_addr; // @[Core.scala 25:19]
  wire [1:0] mmu_io_csr_priv; // @[Core.scala 25:19]
  wire  mmu_io_csr_mxr; // @[Core.scala 25:19]
  wire  mmu_io_csr_sum; // @[Core.scala 25:19]
  wire [31:0] mmu_io_dev_if__addr; // @[Core.scala 25:19]
  wire [3:0] mmu_io_dev_if__mode; // @[Core.scala 25:19]
  wire [31:0] mmu_io_dev_if__rdata; // @[Core.scala 25:19]
  wire  mmu_io_dev_if__ok; // @[Core.scala 25:19]
  wire [31:0] mmu_io_dev_mem_addr; // @[Core.scala 25:19]
  wire [3:0] mmu_io_dev_mem_mode; // @[Core.scala 25:19]
  wire [31:0] mmu_io_dev_mem_wdata; // @[Core.scala 25:19]
  wire [31:0] mmu_io_dev_mem_rdata; // @[Core.scala 25:19]
  wire  mmu_io_dev_mem_ok; // @[Core.scala 25:19]
  wire  csr_clock; // @[Core.scala 26:19]
  wire  csr_reset; // @[Core.scala 26:19]
  wire [11:0] csr_io_id_addr; // @[Core.scala 26:19]
  wire [31:0] csr_io_id_rdata; // @[Core.scala 26:19]
  wire [1:0] csr_io_id_prv; // @[Core.scala 26:19]
  wire  csr_io_mem_wrCSROp_valid; // @[Core.scala 26:19]
  wire [11:0] csr_io_mem_wrCSROp_addr; // @[Core.scala 26:19]
  wire [31:0] csr_io_mem_wrCSROp_data; // @[Core.scala 26:19]
  wire  csr_io_mem_excep_valid; // @[Core.scala 26:19]
  wire [31:0] csr_io_mem_excep_code; // @[Core.scala 26:19]
  wire [31:0] csr_io_mem_excep_value; // @[Core.scala 26:19]
  wire [31:0] csr_io_mem_excep_pc; // @[Core.scala 26:19]
  wire  csr_io_mem_excep_valid_inst; // @[Core.scala 26:19]
  wire  csr_io_mem_inter_valid; // @[Core.scala 26:19]
  wire [31:0] csr_io_mem_inter_bits; // @[Core.scala 26:19]
  wire [31:0] csr_io_mmu_satp; // @[Core.scala 26:19]
  wire  csr_io_mmu_flush_one; // @[Core.scala 26:19]
  wire  csr_io_mmu_flush_all; // @[Core.scala 26:19]
  wire [31:0] csr_io_mmu_flush_addr; // @[Core.scala 26:19]
  wire [1:0] csr_io_mmu_priv; // @[Core.scala 26:19]
  wire  csr_io_mmu_mxr; // @[Core.scala 26:19]
  wire  csr_io_mmu_sum; // @[Core.scala 26:19]
  wire  csr_io_flush; // @[Core.scala 26:19]
  wire [31:0] csr_io_csrNewPc; // @[Core.scala 26:19]
  wire [162:0] _T_10 = {id_io_ex_wrCSROp_data,id_io_ex_store_data,id_io_ex_excep_valid,id_io_ex_excep_code,id_io_ex_excep_value,id_io_ex_excep_pc,id_io_ex_excep_valid_inst,id_io_ex_ready}; // @[Core.scala 63:35]
  wire [282:0] _T_18 = {id_io_ex_aluOp_rd1,id_io_ex_aluOp_rd2,id_io_ex_aluOp_opt,id_io_ex_wrRegOp_addr,33'h0,id_io_ex_wrCSROp_valid,id_io_ex_wrCSROp_addr,_T_10}; // @[Core.scala 63:35]
  IF iff_ ( // @[Core.scala 20:19]
    .clock(iff__clock),
    .reset(iff__reset),
    .io_mmu_addr(iff__io_mmu_addr),
    .io_mmu_mode(iff__io_mmu_mode),
    .io_mmu_rdata(iff__io_mmu_rdata),
    .io_mmu_ok(iff__io_mmu_ok),
    .io_mmu_pageFault(iff__io_mmu_pageFault),
    .io_id_inst(iff__io_id_inst),
    .io_id_excep_valid(iff__io_id_excep_valid),
    .io_id_excep_code(iff__io_id_excep_code),
    .io_id_excep_value(iff__io_id_excep_value),
    .io_id_excep_pc(iff__io_id_excep_pc),
    .io_id_excep_valid_inst(iff__io_id_excep_valid_inst),
    .io_id_branch_valid(iff__io_id_branch_valid),
    .io_id_branch_bits(iff__io_id_branch_bits),
    .io_id_ready(iff__io_id_ready)
  );
  ID id ( // @[Core.scala 21:19]
    .clock(id_clock),
    .reset(id_reset),
    .io_iff_inst(id_io_iff_inst),
    .io_iff_excep_valid(id_io_iff_excep_valid),
    .io_iff_excep_code(id_io_iff_excep_code),
    .io_iff_excep_value(id_io_iff_excep_value),
    .io_iff_excep_pc(id_io_iff_excep_pc),
    .io_iff_excep_valid_inst(id_io_iff_excep_valid_inst),
    .io_iff_branch_valid(id_io_iff_branch_valid),
    .io_iff_branch_bits(id_io_iff_branch_bits),
    .io_iff_ready(id_io_iff_ready),
    .io_reg_read1_addr(id_io_reg_read1_addr),
    .io_reg_read1_data(id_io_reg_read1_data),
    .io_reg_read2_addr(id_io_reg_read2_addr),
    .io_reg_read2_data(id_io_reg_read2_data),
    .io_ex_aluOp_rd1(id_io_ex_aluOp_rd1),
    .io_ex_aluOp_rd2(id_io_ex_aluOp_rd2),
    .io_ex_aluOp_opt(id_io_ex_aluOp_opt),
    .io_ex_wrRegOp_addr(id_io_ex_wrRegOp_addr),
    .io_ex_wrCSROp_valid(id_io_ex_wrCSROp_valid),
    .io_ex_wrCSROp_addr(id_io_ex_wrCSROp_addr),
    .io_ex_wrCSROp_data(id_io_ex_wrCSROp_data),
    .io_ex_store_data(id_io_ex_store_data),
    .io_ex_excep_valid(id_io_ex_excep_valid),
    .io_ex_excep_code(id_io_ex_excep_code),
    .io_ex_excep_value(id_io_ex_excep_value),
    .io_ex_excep_pc(id_io_ex_excep_pc),
    .io_ex_excep_valid_inst(id_io_ex_excep_valid_inst),
    .io_ex_ready(id_io_ex_ready),
    .io_csr_addr(id_io_csr_addr),
    .io_csr_rdata(id_io_csr_rdata),
    .io_csr_prv(id_io_csr_prv),
    .io_flush(id_io_flush),
    .io_exWrRegOp_addr(id_io_exWrRegOp_addr),
    .io_exWrRegOp_data(id_io_exWrRegOp_data),
    .io_exWrRegOp_rdy(id_io_exWrRegOp_rdy),
    .io_memWrRegOp_addr(id_io_memWrRegOp_addr),
    .io_memWrRegOp_data(id_io_memWrRegOp_data),
    .io_exWrCSROp_valid(id_io_exWrCSROp_valid),
    .io_exWrCSROp_addr(id_io_exWrCSROp_addr),
    .io_exWrCSROp_data(id_io_exWrCSROp_data),
    .io_memWrCSROp_valid(id_io_memWrCSROp_valid),
    .io_memWrCSROp_addr(id_io_memWrCSROp_addr),
    .io_memWrCSROp_data(id_io_memWrCSROp_data)
  );
  EX ex ( // @[Core.scala 22:19]
    .clock(ex_clock),
    .reset(ex_reset),
    .io_id_aluOp_rd1(ex_io_id_aluOp_rd1),
    .io_id_aluOp_rd2(ex_io_id_aluOp_rd2),
    .io_id_aluOp_opt(ex_io_id_aluOp_opt),
    .io_id_wrRegOp_addr(ex_io_id_wrRegOp_addr),
    .io_id_wrCSROp_valid(ex_io_id_wrCSROp_valid),
    .io_id_wrCSROp_addr(ex_io_id_wrCSROp_addr),
    .io_id_wrCSROp_data(ex_io_id_wrCSROp_data),
    .io_id_store_data(ex_io_id_store_data),
    .io_id_excep_valid(ex_io_id_excep_valid),
    .io_id_excep_code(ex_io_id_excep_code),
    .io_id_excep_value(ex_io_id_excep_value),
    .io_id_excep_pc(ex_io_id_excep_pc),
    .io_id_excep_valid_inst(ex_io_id_excep_valid_inst),
    .io_id_ready(ex_io_id_ready),
    .io_mem_ramOp_addr(ex_io_mem_ramOp_addr),
    .io_mem_ramOp_mode(ex_io_mem_ramOp_mode),
    .io_mem_ramOp_wdata(ex_io_mem_ramOp_wdata),
    .io_mem_wrRegOp_addr(ex_io_mem_wrRegOp_addr),
    .io_mem_wrRegOp_data(ex_io_mem_wrRegOp_data),
    .io_mem_wrRegOp_rdy(ex_io_mem_wrRegOp_rdy),
    .io_mem_wrCSROp_valid(ex_io_mem_wrCSROp_valid),
    .io_mem_wrCSROp_addr(ex_io_mem_wrCSROp_addr),
    .io_mem_wrCSROp_data(ex_io_mem_wrCSROp_data),
    .io_mem_excep_valid(ex_io_mem_excep_valid),
    .io_mem_excep_code(ex_io_mem_excep_code),
    .io_mem_excep_value(ex_io_mem_excep_value),
    .io_mem_excep_pc(ex_io_mem_excep_pc),
    .io_mem_excep_valid_inst(ex_io_mem_excep_valid_inst),
    .io_mem_ready(ex_io_mem_ready),
    .io_flush(ex_io_flush)
  );
  MEM mem ( // @[Core.scala 23:19]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_ex_ramOp_addr(mem_io_ex_ramOp_addr),
    .io_ex_ramOp_mode(mem_io_ex_ramOp_mode),
    .io_ex_ramOp_wdata(mem_io_ex_ramOp_wdata),
    .io_ex_wrRegOp_addr(mem_io_ex_wrRegOp_addr),
    .io_ex_wrRegOp_data(mem_io_ex_wrRegOp_data),
    .io_ex_wrCSROp_valid(mem_io_ex_wrCSROp_valid),
    .io_ex_wrCSROp_addr(mem_io_ex_wrCSROp_addr),
    .io_ex_wrCSROp_data(mem_io_ex_wrCSROp_data),
    .io_ex_excep_valid(mem_io_ex_excep_valid),
    .io_ex_excep_code(mem_io_ex_excep_code),
    .io_ex_excep_value(mem_io_ex_excep_value),
    .io_ex_excep_pc(mem_io_ex_excep_pc),
    .io_ex_excep_valid_inst(mem_io_ex_excep_valid_inst),
    .io_ex_ready(mem_io_ex_ready),
    .io_mmu_addr(mem_io_mmu_addr),
    .io_mmu_mode(mem_io_mmu_mode),
    .io_mmu_wdata(mem_io_mmu_wdata),
    .io_mmu_rdata(mem_io_mmu_rdata),
    .io_mmu_ok(mem_io_mmu_ok),
    .io_mmu_pageFault(mem_io_mmu_pageFault),
    .io_csr_wrCSROp_valid(mem_io_csr_wrCSROp_valid),
    .io_csr_wrCSROp_addr(mem_io_csr_wrCSROp_addr),
    .io_csr_wrCSROp_data(mem_io_csr_wrCSROp_data),
    .io_csr_excep_valid(mem_io_csr_excep_valid),
    .io_csr_excep_code(mem_io_csr_excep_code),
    .io_csr_excep_value(mem_io_csr_excep_value),
    .io_csr_excep_pc(mem_io_csr_excep_pc),
    .io_csr_excep_valid_inst(mem_io_csr_excep_valid_inst),
    .io_csr_inter_valid(mem_io_csr_inter_valid),
    .io_csr_inter_bits(mem_io_csr_inter_bits),
    .io_reg_addr(mem_io_reg_addr),
    .io_reg_data(mem_io_reg_data),
    .io_flush(mem_io_flush)
  );
  RegFile reg_ ( // @[Core.scala 24:19]
    .clock(reg__clock),
    .io_id_read1_addr(reg__io_id_read1_addr),
    .io_id_read1_data(reg__io_id_read1_data),
    .io_id_read2_addr(reg__io_id_read2_addr),
    .io_id_read2_data(reg__io_id_read2_data),
    .io_mem_addr(reg__io_mem_addr),
    .io_mem_data(reg__io_mem_data),
    .io_log_0(reg__io_log_0),
    .io_log_1(reg__io_log_1),
    .io_log_2(reg__io_log_2),
    .io_log_3(reg__io_log_3),
    .io_log_4(reg__io_log_4),
    .io_log_5(reg__io_log_5),
    .io_log_6(reg__io_log_6),
    .io_log_7(reg__io_log_7),
    .io_log_8(reg__io_log_8),
    .io_log_9(reg__io_log_9),
    .io_log_10(reg__io_log_10),
    .io_log_11(reg__io_log_11),
    .io_log_12(reg__io_log_12),
    .io_log_13(reg__io_log_13),
    .io_log_14(reg__io_log_14),
    .io_log_15(reg__io_log_15),
    .io_log_16(reg__io_log_16),
    .io_log_17(reg__io_log_17),
    .io_log_18(reg__io_log_18),
    .io_log_19(reg__io_log_19),
    .io_log_20(reg__io_log_20),
    .io_log_21(reg__io_log_21),
    .io_log_22(reg__io_log_22),
    .io_log_23(reg__io_log_23),
    .io_log_24(reg__io_log_24),
    .io_log_25(reg__io_log_25),
    .io_log_26(reg__io_log_26),
    .io_log_27(reg__io_log_27),
    .io_log_28(reg__io_log_28),
    .io_log_29(reg__io_log_29),
    .io_log_30(reg__io_log_30),
    .io_log_31(reg__io_log_31)
  );
  MMU mmu ( // @[Core.scala 25:19]
    .clock(mmu_clock),
    .reset(mmu_reset),
    .io_iff_addr(mmu_io_iff_addr),
    .io_iff_mode(mmu_io_iff_mode),
    .io_iff_rdata(mmu_io_iff_rdata),
    .io_iff_ok(mmu_io_iff_ok),
    .io_iff_pageFault(mmu_io_iff_pageFault),
    .io_mem_addr(mmu_io_mem_addr),
    .io_mem_mode(mmu_io_mem_mode),
    .io_mem_wdata(mmu_io_mem_wdata),
    .io_mem_rdata(mmu_io_mem_rdata),
    .io_mem_ok(mmu_io_mem_ok),
    .io_mem_pageFault(mmu_io_mem_pageFault),
    .io_csr_satp(mmu_io_csr_satp),
    .io_csr_flush_one(mmu_io_csr_flush_one),
    .io_csr_flush_all(mmu_io_csr_flush_all),
    .io_csr_flush_addr(mmu_io_csr_flush_addr),
    .io_csr_priv(mmu_io_csr_priv),
    .io_csr_mxr(mmu_io_csr_mxr),
    .io_csr_sum(mmu_io_csr_sum),
    .io_dev_if__addr(mmu_io_dev_if__addr),
    .io_dev_if__mode(mmu_io_dev_if__mode),
    .io_dev_if__rdata(mmu_io_dev_if__rdata),
    .io_dev_if__ok(mmu_io_dev_if__ok),
    .io_dev_mem_addr(mmu_io_dev_mem_addr),
    .io_dev_mem_mode(mmu_io_dev_mem_mode),
    .io_dev_mem_wdata(mmu_io_dev_mem_wdata),
    .io_dev_mem_rdata(mmu_io_dev_mem_rdata),
    .io_dev_mem_ok(mmu_io_dev_mem_ok)
  );
  CSR csr ( // @[Core.scala 26:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_id_addr(csr_io_id_addr),
    .io_id_rdata(csr_io_id_rdata),
    .io_id_prv(csr_io_id_prv),
    .io_mem_wrCSROp_valid(csr_io_mem_wrCSROp_valid),
    .io_mem_wrCSROp_addr(csr_io_mem_wrCSROp_addr),
    .io_mem_wrCSROp_data(csr_io_mem_wrCSROp_data),
    .io_mem_excep_valid(csr_io_mem_excep_valid),
    .io_mem_excep_code(csr_io_mem_excep_code),
    .io_mem_excep_value(csr_io_mem_excep_value),
    .io_mem_excep_pc(csr_io_mem_excep_pc),
    .io_mem_excep_valid_inst(csr_io_mem_excep_valid_inst),
    .io_mem_inter_valid(csr_io_mem_inter_valid),
    .io_mem_inter_bits(csr_io_mem_inter_bits),
    .io_mmu_satp(csr_io_mmu_satp),
    .io_mmu_flush_one(csr_io_mmu_flush_one),
    .io_mmu_flush_all(csr_io_mmu_flush_all),
    .io_mmu_flush_addr(csr_io_mmu_flush_addr),
    .io_mmu_priv(csr_io_mmu_priv),
    .io_mmu_mxr(csr_io_mmu_mxr),
    .io_mmu_sum(csr_io_mmu_sum),
    .io_flush(csr_io_flush),
    .io_csrNewPc(csr_io_csrNewPc)
  );
  assign io_dev_if__addr = mmu_io_dev_if__addr; // @[Core.scala 46:20]
  assign io_dev_if__mode = mmu_io_dev_if__mode; // @[Core.scala 46:20]
  assign io_dev_mem_addr = mmu_io_dev_mem_addr; // @[Core.scala 46:20]
  assign io_dev_mem_mode = mmu_io_dev_mem_mode; // @[Core.scala 46:20]
  assign io_dev_mem_wdata = mmu_io_dev_mem_wdata; // @[Core.scala 46:20]
  assign io_debug_idex_aluOp_rd1 = _T_18[281:250]; // @[Core.scala 63:15]
  assign io_debug_idex_aluOp_rd2 = _T_18[249:218]; // @[Core.scala 63:15]
  assign io_debug_idex_aluOp_opt = _T_18[217:213]; // @[Core.scala 63:15]
  assign io_debug_idex_wrRegOp_addr = _T_18[212:208]; // @[Core.scala 63:15]
  assign io_debug_idex_wrRegOp_data = _T_18[207:176]; // @[Core.scala 63:15]
  assign io_debug_idex_wrRegOp_rdy = _T_18[175]; // @[Core.scala 63:15]
  assign io_debug_idex_wrCSROp_valid = _T_18[174]; // @[Core.scala 63:15]
  assign io_debug_idex_wrCSROp_addr = _T_18[173:162]; // @[Core.scala 63:15]
  assign io_debug_idex_wrCSROp_data = _T_18[161:130]; // @[Core.scala 63:15]
  assign io_debug_idex_store_data = _T_18[129:98]; // @[Core.scala 63:15]
  assign io_debug_idex_excep_valid = _T_18[97]; // @[Core.scala 63:15]
  assign io_debug_idex_excep_code = _T_18[96:65]; // @[Core.scala 63:15]
  assign io_debug_idex_excep_value = _T_18[64:33]; // @[Core.scala 63:15]
  assign io_debug_idex_excep_pc = _T_18[32:1]; // @[Core.scala 63:15]
  assign io_debug_idex_excep_valid_inst = _T_18[0]; // @[Core.scala 63:15]
  assign io_debug_ifpc = iff__io_id_excep_pc; // @[Core.scala 62:15]
  assign io_debug_reg_0 = reg__io_log_0; // @[Core.scala 61:15]
  assign io_debug_reg_1 = reg__io_log_1; // @[Core.scala 61:15]
  assign io_debug_reg_2 = reg__io_log_2; // @[Core.scala 61:15]
  assign io_debug_reg_3 = reg__io_log_3; // @[Core.scala 61:15]
  assign io_debug_reg_4 = reg__io_log_4; // @[Core.scala 61:15]
  assign io_debug_reg_5 = reg__io_log_5; // @[Core.scala 61:15]
  assign io_debug_reg_6 = reg__io_log_6; // @[Core.scala 61:15]
  assign io_debug_reg_7 = reg__io_log_7; // @[Core.scala 61:15]
  assign io_debug_reg_8 = reg__io_log_8; // @[Core.scala 61:15]
  assign io_debug_reg_9 = reg__io_log_9; // @[Core.scala 61:15]
  assign io_debug_reg_10 = reg__io_log_10; // @[Core.scala 61:15]
  assign io_debug_reg_11 = reg__io_log_11; // @[Core.scala 61:15]
  assign io_debug_reg_12 = reg__io_log_12; // @[Core.scala 61:15]
  assign io_debug_reg_13 = reg__io_log_13; // @[Core.scala 61:15]
  assign io_debug_reg_14 = reg__io_log_14; // @[Core.scala 61:15]
  assign io_debug_reg_15 = reg__io_log_15; // @[Core.scala 61:15]
  assign io_debug_reg_16 = reg__io_log_16; // @[Core.scala 61:15]
  assign io_debug_reg_17 = reg__io_log_17; // @[Core.scala 61:15]
  assign io_debug_reg_18 = reg__io_log_18; // @[Core.scala 61:15]
  assign io_debug_reg_19 = reg__io_log_19; // @[Core.scala 61:15]
  assign io_debug_reg_20 = reg__io_log_20; // @[Core.scala 61:15]
  assign io_debug_reg_21 = reg__io_log_21; // @[Core.scala 61:15]
  assign io_debug_reg_22 = reg__io_log_22; // @[Core.scala 61:15]
  assign io_debug_reg_23 = reg__io_log_23; // @[Core.scala 61:15]
  assign io_debug_reg_24 = reg__io_log_24; // @[Core.scala 61:15]
  assign io_debug_reg_25 = reg__io_log_25; // @[Core.scala 61:15]
  assign io_debug_reg_26 = reg__io_log_26; // @[Core.scala 61:15]
  assign io_debug_reg_27 = reg__io_log_27; // @[Core.scala 61:15]
  assign io_debug_reg_28 = reg__io_log_28; // @[Core.scala 61:15]
  assign io_debug_reg_29 = reg__io_log_29; // @[Core.scala 61:15]
  assign io_debug_reg_30 = reg__io_log_30; // @[Core.scala 61:15]
  assign io_debug_reg_31 = reg__io_log_31; // @[Core.scala 61:15]
  assign io_debug_finish_pc_valid = mem_io_csr_excep_valid_inst; // @[Core.scala 64:21]
  assign io_debug_finish_pc_bits = mem_io_csr_excep_pc; // @[Core.scala 65:21]
  assign iff__clock = clock;
  assign iff__reset = reset;
  assign iff__io_mmu_rdata = mmu_io_iff_rdata; // @[Core.scala 44:20]
  assign iff__io_mmu_ok = mmu_io_iff_ok; // @[Core.scala 44:20]
  assign iff__io_mmu_pageFault = mmu_io_iff_pageFault; // @[Core.scala 44:20]
  assign iff__io_id_branch_valid = csr_io_flush | id_io_iff_branch_valid; // @[Core.scala 29:20 Core.scala 50:26]
  assign iff__io_id_branch_bits = csr_io_flush ? csr_io_csrNewPc : id_io_iff_branch_bits; // @[Core.scala 29:20 Core.scala 51:25]
  assign iff__io_id_ready = id_io_iff_ready; // @[Core.scala 29:20]
  assign id_clock = clock;
  assign id_reset = reset;
  assign id_io_iff_inst = iff__io_id_inst; // @[Core.scala 29:20]
  assign id_io_iff_excep_valid = iff__io_id_excep_valid; // @[Core.scala 29:20]
  assign id_io_iff_excep_code = iff__io_id_excep_code; // @[Core.scala 29:20]
  assign id_io_iff_excep_value = iff__io_id_excep_value; // @[Core.scala 29:20]
  assign id_io_iff_excep_pc = iff__io_id_excep_pc; // @[Core.scala 29:20]
  assign id_io_iff_excep_valid_inst = iff__io_id_excep_valid_inst; // @[Core.scala 29:20]
  assign id_io_reg_read1_data = reg__io_id_read1_data; // @[Core.scala 36:20]
  assign id_io_reg_read2_data = reg__io_id_read2_data; // @[Core.scala 36:20]
  assign id_io_ex_ready = ex_io_id_ready; // @[Core.scala 30:20]
  assign id_io_csr_rdata = csr_io_id_rdata; // @[Core.scala 37:20]
  assign id_io_csr_prv = csr_io_id_prv; // @[Core.scala 37:20]
  assign id_io_flush = csr_io_flush; // @[Core.scala 52:15]
  assign id_io_exWrRegOp_addr = ex_io_mem_wrRegOp_addr; // @[Core.scala 38:20]
  assign id_io_exWrRegOp_data = ex_io_mem_wrRegOp_data; // @[Core.scala 38:20]
  assign id_io_exWrRegOp_rdy = ex_io_mem_wrRegOp_rdy; // @[Core.scala 38:20]
  assign id_io_memWrRegOp_addr = mem_io_reg_addr; // @[Core.scala 39:20]
  assign id_io_memWrRegOp_data = mem_io_reg_data; // @[Core.scala 39:20]
  assign id_io_exWrCSROp_valid = ex_io_mem_wrCSROp_valid; // @[Core.scala 40:20]
  assign id_io_exWrCSROp_addr = ex_io_mem_wrCSROp_addr; // @[Core.scala 40:20]
  assign id_io_exWrCSROp_data = ex_io_mem_wrCSROp_data; // @[Core.scala 40:20]
  assign id_io_memWrCSROp_valid = mem_io_csr_wrCSROp_valid; // @[Core.scala 41:20]
  assign id_io_memWrCSROp_addr = mem_io_csr_wrCSROp_addr; // @[Core.scala 41:20]
  assign id_io_memWrCSROp_data = mem_io_csr_wrCSROp_data; // @[Core.scala 41:20]
  assign ex_clock = clock;
  assign ex_reset = reset;
  assign ex_io_id_aluOp_rd1 = id_io_ex_aluOp_rd1; // @[Core.scala 30:20]
  assign ex_io_id_aluOp_rd2 = id_io_ex_aluOp_rd2; // @[Core.scala 30:20]
  assign ex_io_id_aluOp_opt = id_io_ex_aluOp_opt; // @[Core.scala 30:20]
  assign ex_io_id_wrRegOp_addr = id_io_ex_wrRegOp_addr; // @[Core.scala 30:20]
  assign ex_io_id_wrCSROp_valid = id_io_ex_wrCSROp_valid; // @[Core.scala 30:20]
  assign ex_io_id_wrCSROp_addr = id_io_ex_wrCSROp_addr; // @[Core.scala 30:20]
  assign ex_io_id_wrCSROp_data = id_io_ex_wrCSROp_data; // @[Core.scala 30:20]
  assign ex_io_id_store_data = id_io_ex_store_data; // @[Core.scala 30:20]
  assign ex_io_id_excep_valid = id_io_ex_excep_valid; // @[Core.scala 30:20]
  assign ex_io_id_excep_code = id_io_ex_excep_code; // @[Core.scala 30:20]
  assign ex_io_id_excep_value = id_io_ex_excep_value; // @[Core.scala 30:20]
  assign ex_io_id_excep_pc = id_io_ex_excep_pc; // @[Core.scala 30:20]
  assign ex_io_id_excep_valid_inst = id_io_ex_excep_valid_inst; // @[Core.scala 30:20]
  assign ex_io_mem_ready = mem_io_ex_ready; // @[Core.scala 31:20]
  assign ex_io_flush = csr_io_flush; // @[Core.scala 53:15]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_ex_ramOp_addr = ex_io_mem_ramOp_addr; // @[Core.scala 31:20]
  assign mem_io_ex_ramOp_mode = ex_io_mem_ramOp_mode; // @[Core.scala 31:20]
  assign mem_io_ex_ramOp_wdata = ex_io_mem_ramOp_wdata; // @[Core.scala 31:20]
  assign mem_io_ex_wrRegOp_addr = ex_io_mem_wrRegOp_addr; // @[Core.scala 31:20]
  assign mem_io_ex_wrRegOp_data = ex_io_mem_wrRegOp_data; // @[Core.scala 31:20]
  assign mem_io_ex_wrCSROp_valid = ex_io_mem_wrCSROp_valid; // @[Core.scala 31:20]
  assign mem_io_ex_wrCSROp_addr = ex_io_mem_wrCSROp_addr; // @[Core.scala 31:20]
  assign mem_io_ex_wrCSROp_data = ex_io_mem_wrCSROp_data; // @[Core.scala 31:20]
  assign mem_io_ex_excep_valid = ex_io_mem_excep_valid; // @[Core.scala 31:20]
  assign mem_io_ex_excep_code = ex_io_mem_excep_code; // @[Core.scala 31:20]
  assign mem_io_ex_excep_value = ex_io_mem_excep_value; // @[Core.scala 31:20]
  assign mem_io_ex_excep_pc = ex_io_mem_excep_pc; // @[Core.scala 31:20]
  assign mem_io_ex_excep_valid_inst = ex_io_mem_excep_valid_inst; // @[Core.scala 31:20]
  assign mem_io_mmu_rdata = mmu_io_mem_rdata; // @[Core.scala 45:20]
  assign mem_io_mmu_ok = mmu_io_mem_ok; // @[Core.scala 45:20]
  assign mem_io_mmu_pageFault = mmu_io_mem_pageFault; // @[Core.scala 45:20]
  assign mem_io_csr_inter_valid = csr_io_mem_inter_valid; // @[Core.scala 33:20]
  assign mem_io_csr_inter_bits = csr_io_mem_inter_bits; // @[Core.scala 33:20]
  assign mem_io_flush = csr_io_flush; // @[Core.scala 54:16]
  assign reg__clock = clock;
  assign reg__io_id_read1_addr = id_io_reg_read1_addr; // @[Core.scala 36:20]
  assign reg__io_id_read2_addr = id_io_reg_read2_addr; // @[Core.scala 36:20]
  assign reg__io_mem_addr = mem_io_reg_addr; // @[Core.scala 32:20]
  assign reg__io_mem_data = mem_io_reg_data; // @[Core.scala 32:20]
  assign mmu_clock = clock;
  assign mmu_reset = reset;
  assign mmu_io_iff_addr = iff__io_mmu_addr; // @[Core.scala 44:20]
  assign mmu_io_iff_mode = iff__io_mmu_mode; // @[Core.scala 44:20]
  assign mmu_io_mem_addr = mem_io_mmu_addr; // @[Core.scala 45:20]
  assign mmu_io_mem_mode = mem_io_mmu_mode; // @[Core.scala 45:20]
  assign mmu_io_mem_wdata = mem_io_mmu_wdata; // @[Core.scala 45:20]
  assign mmu_io_csr_satp = csr_io_mmu_satp; // @[Core.scala 47:20]
  assign mmu_io_csr_flush_one = csr_io_mmu_flush_one; // @[Core.scala 47:20]
  assign mmu_io_csr_flush_all = csr_io_mmu_flush_all; // @[Core.scala 47:20]
  assign mmu_io_csr_flush_addr = csr_io_mmu_flush_addr; // @[Core.scala 47:20]
  assign mmu_io_csr_priv = csr_io_mmu_priv; // @[Core.scala 47:20]
  assign mmu_io_csr_mxr = csr_io_mmu_mxr; // @[Core.scala 47:20]
  assign mmu_io_csr_sum = csr_io_mmu_sum; // @[Core.scala 47:20]
  assign mmu_io_dev_if__rdata = io_dev_if__rdata; // @[Core.scala 46:20]
  assign mmu_io_dev_if__ok = io_dev_if__ok; // @[Core.scala 46:20]
  assign mmu_io_dev_mem_rdata = io_dev_mem_rdata; // @[Core.scala 46:20]
  assign mmu_io_dev_mem_ok = io_dev_mem_ok; // @[Core.scala 46:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_id_addr = id_io_csr_addr; // @[Core.scala 37:20]
  assign csr_io_mem_wrCSROp_valid = mem_io_csr_wrCSROp_valid; // @[Core.scala 33:20]
  assign csr_io_mem_wrCSROp_addr = mem_io_csr_wrCSROp_addr; // @[Core.scala 33:20]
  assign csr_io_mem_wrCSROp_data = mem_io_csr_wrCSROp_data; // @[Core.scala 33:20]
  assign csr_io_mem_excep_valid = mem_io_csr_excep_valid; // @[Core.scala 33:20]
  assign csr_io_mem_excep_code = mem_io_csr_excep_code; // @[Core.scala 33:20]
  assign csr_io_mem_excep_value = mem_io_csr_excep_value; // @[Core.scala 33:20]
  assign csr_io_mem_excep_pc = mem_io_csr_excep_pc; // @[Core.scala 33:20]
  assign csr_io_mem_excep_valid_inst = mem_io_csr_excep_valid_inst; // @[Core.scala 33:20]
endmodule
module IOManager(
  input         clock,
  input         reset,
  input  [31:0] io_core_if__addr,
  input  [3:0]  io_core_if__mode,
  output [31:0] io_core_if__rdata,
  output        io_core_if__ok,
  input  [31:0] io_core_mem_addr,
  input  [3:0]  io_core_mem_mode,
  input  [31:0] io_core_mem_wdata,
  output [31:0] io_core_mem_rdata,
  output        io_core_mem_ok,
  output [31:0] io_ram_addr,
  output [3:0]  io_ram_mode,
  output [31:0] io_ram_wdata,
  input  [31:0] io_ram_rdata,
  input         io_ram_ok,
  output [31:0] io_flash_addr,
  output [3:0]  io_flash_mode,
  output [31:0] io_flash_wdata,
  input  [31:0] io_flash_rdata,
  input         io_flash_ok,
  output [31:0] io_serial_addr,
  output [3:0]  io_serial_mode,
  output [31:0] io_serial_wdata,
  input  [31:0] io_serial_rdata,
  input         io_serial_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ifWait; // @[IOManager.scala 69:24]
  reg [1:0] memWait; // @[IOManager.scala 70:24]
  wire  _T = 2'h1 == ifWait; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h2 == ifWait; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h3 == ifWait; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_0 = _T_2 ? io_serial_rdata : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_1 = _T_2 & io_serial_ok; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_2 = _T_1 ? io_flash_rdata : _GEN_0; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_1 ? io_flash_ok : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T ? io_ram_ok : _GEN_3; // @[Conditional.scala 40:58]
  wire  _T_3 = 2'h1 == memWait; // @[Conditional.scala 37:30]
  wire  _T_4 = 2'h2 == memWait; // @[Conditional.scala 37:30]
  wire  _T_5 = 2'h3 == memWait; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_6 = _T_5 ? io_serial_rdata : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_5 & io_serial_ok; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_8 = _T_4 ? io_flash_rdata : _GEN_6; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_4 ? io_flash_ok : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_3 ? io_ram_ok : _GEN_9; // @[Conditional.scala 40:58]
  wire  _T_6 = ifWait != 2'h2; // @[IOManager.scala 93:26]
  wire  _T_7 = memWait != 2'h2; // @[IOManager.scala 93:51]
  wire  flashFree = _T_6 & _T_7; // @[IOManager.scala 93:40]
  wire  _T_8 = ifWait != 2'h0; // @[IOManager.scala 94:24]
  wire  _T_9 = ~io_core_if__ok; // @[IOManager.scala 94:40]
  wire  _T_10 = _T_8 & _T_9; // @[IOManager.scala 94:37]
  wire  _T_12 = memWait != 2'h0; // @[IOManager.scala 95:26]
  wire  _T_13 = ~io_core_mem_ok; // @[IOManager.scala 95:42]
  wire  _T_14 = _T_12 & _T_13; // @[IOManager.scala 95:39]
  wire  _T_16 = memWait == 2'h0; // @[IOManager.scala 98:16]
  wire  _T_17 = io_core_mem_mode != 4'h0; // @[IOManager.scala 98:41]
  wire  _T_18 = _T_16 & _T_17; // @[IOManager.scala 98:29]
  wire  _T_19 = io_core_mem_addr >= 32'h80000000; // @[IOManager.scala 16:22]
  wire  _T_20 = io_core_mem_addr < 32'h80800000; // @[IOManager.scala 16:43]
  wire  _T_21 = _T_19 & _T_20; // @[IOManager.scala 16:35]
  wire  _T_23 = io_core_mem_addr >= 32'h800000; // @[IOManager.scala 17:24]
  wire  _T_24 = io_core_mem_addr < 32'h1000000; // @[IOManager.scala 17:47]
  wire  _T_25 = _T_23 & _T_24; // @[IOManager.scala 17:39]
  wire [3:0] _GEN_14 = flashFree ? io_core_mem_mode : 4'h0; // @[IOManager.scala 109:23]
  wire [31:0] _GEN_15 = flashFree ? io_core_mem_addr : 32'h0; // @[IOManager.scala 109:23]
  wire [31:0] _GEN_16 = flashFree ? io_core_mem_wdata : 32'h0; // @[IOManager.scala 109:23]
  wire  _T_26 = io_core_mem_addr >= 32'h10000000; // @[IOManager.scala 18:25]
  wire  _T_27 = io_core_mem_addr < 32'h10000008; // @[IOManager.scala 18:49]
  wire  _T_28 = _T_26 & _T_27; // @[IOManager.scala 18:41]
  wire  _T_31 = ~reset; // @[IOManager.scala 123:13]
  wire [3:0] _GEN_20 = _T_28 ? io_core_mem_mode : 4'h0; // @[IOManager.scala 113:35]
  wire [31:0] _GEN_21 = _T_28 ? io_core_mem_addr : 32'h0; // @[IOManager.scala 113:35]
  wire [31:0] _GEN_22 = _T_28 ? io_core_mem_wdata : 32'h0; // @[IOManager.scala 113:35]
  wire  _GEN_24 = _T_28 ? io_core_mem_mode[3] : _GEN_11; // @[IOManager.scala 113:35]
  wire [3:0] _GEN_25 = _T_25 ? _GEN_14 : 4'h0; // @[IOManager.scala 108:34]
  wire [31:0] _GEN_26 = _T_25 ? _GEN_15 : 32'h0; // @[IOManager.scala 108:34]
  wire [31:0] _GEN_27 = _T_25 ? _GEN_16 : 32'h0; // @[IOManager.scala 108:34]
  wire [3:0] _GEN_29 = _T_25 ? 4'h0 : _GEN_20; // @[IOManager.scala 108:34]
  wire [31:0] _GEN_30 = _T_25 ? 32'h0 : _GEN_21; // @[IOManager.scala 108:34]
  wire [31:0] _GEN_31 = _T_25 ? 32'h0 : _GEN_22; // @[IOManager.scala 108:34]
  wire  _GEN_32 = _T_25 ? _GEN_11 : _GEN_24; // @[IOManager.scala 108:34]
  wire [3:0] _GEN_33 = _T_21 ? io_core_mem_mode : 4'h0; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_34 = _T_21 ? io_core_mem_addr : 32'h0; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_35 = _T_21 ? io_core_mem_wdata : 32'h0; // @[IOManager.scala 99:26]
  wire  _GEN_37 = _T_21 ? io_core_mem_mode[3] : _GEN_32; // @[IOManager.scala 99:26]
  wire [3:0] _GEN_38 = _T_21 ? 4'h0 : _GEN_25; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_39 = _T_21 ? 32'h0 : _GEN_26; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_40 = _T_21 ? 32'h0 : _GEN_27; // @[IOManager.scala 99:26]
  wire [3:0] _GEN_41 = _T_21 ? 4'h0 : _GEN_29; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_42 = _T_21 ? 32'h0 : _GEN_30; // @[IOManager.scala 99:26]
  wire [31:0] _GEN_43 = _T_21 ? 32'h0 : _GEN_31; // @[IOManager.scala 99:26]
  wire [3:0] _GEN_44 = _T_18 ? _GEN_33 : 4'h0; // @[IOManager.scala 98:58]
  wire [31:0] _GEN_45 = _T_18 ? _GEN_34 : 32'h0; // @[IOManager.scala 98:58]
  wire [31:0] _GEN_46 = _T_18 ? _GEN_35 : 32'h0; // @[IOManager.scala 98:58]
  wire [3:0] _GEN_49 = _T_18 ? _GEN_38 : 4'h0; // @[IOManager.scala 98:58]
  wire [31:0] _GEN_50 = _T_18 ? _GEN_39 : 32'h0; // @[IOManager.scala 98:58]
  wire [31:0] _GEN_51 = _T_18 ? _GEN_40 : 32'h0; // @[IOManager.scala 98:58]
  wire  _T_32 = ifWait == 2'h0; // @[IOManager.scala 129:15]
  wire  _T_34 = _T_32 & _T_16; // @[IOManager.scala 129:28]
  wire  _T_35 = io_core_mem_mode == 4'h0; // @[IOManager.scala 129:64]
  wire  _T_36 = _T_34 & _T_35; // @[IOManager.scala 129:52]
  wire  _T_37 = io_core_if__mode != 4'h0; // @[IOManager.scala 129:92]
  wire  _T_38 = _T_36 & _T_37; // @[IOManager.scala 129:80]
  wire  _T_39 = io_core_if__addr >= 32'h80000000; // @[IOManager.scala 16:22]
  wire  _T_40 = io_core_if__addr < 32'h80800000; // @[IOManager.scala 16:43]
  wire  _T_41 = _T_39 & _T_40; // @[IOManager.scala 16:35]
  wire  _T_42 = io_core_if__addr >= 32'h800000; // @[IOManager.scala 17:24]
  wire  _T_43 = io_core_if__addr < 32'h1000000; // @[IOManager.scala 17:47]
  wire  _T_44 = _T_42 & _T_43; // @[IOManager.scala 17:39]
  wire [3:0] _GEN_55 = _T_44 ? io_core_if__mode : _GEN_49; // @[IOManager.scala 134:34]
  wire [31:0] _GEN_56 = _T_44 ? io_core_if__addr : _GEN_50; // @[IOManager.scala 134:34]
  wire [31:0] _GEN_57 = _T_44 ? 32'h0 : _GEN_51; // @[IOManager.scala 134:34]
  wire  _GEN_59 = _T_44 ? 1'h0 : _GEN_5; // @[IOManager.scala 134:34]
  wire [3:0] _GEN_60 = _T_41 ? io_core_if__mode : _GEN_44; // @[IOManager.scala 130:26]
  wire [31:0] _GEN_61 = _T_41 ? io_core_if__addr : _GEN_45; // @[IOManager.scala 130:26]
  wire [31:0] _GEN_62 = _T_41 ? 32'h0 : _GEN_46; // @[IOManager.scala 130:26]
  wire  _GEN_64 = _T_41 ? 1'h0 : _GEN_59; // @[IOManager.scala 130:26]
  wire [3:0] _GEN_65 = _T_41 ? _GEN_49 : _GEN_55; // @[IOManager.scala 130:26]
  wire [31:0] _GEN_66 = _T_41 ? _GEN_50 : _GEN_56; // @[IOManager.scala 130:26]
  wire [31:0] _GEN_67 = _T_41 ? _GEN_51 : _GEN_57; // @[IOManager.scala 130:26]
  wire  _GEN_76 = ~_T_21; // @[IOManager.scala 123:13]
  wire  _GEN_77 = _T_18 & _GEN_76; // @[IOManager.scala 123:13]
  wire  _GEN_78 = ~_T_25; // @[IOManager.scala 123:13]
  wire  _GEN_79 = _GEN_77 & _GEN_78; // @[IOManager.scala 123:13]
  wire  _GEN_80 = ~_T_28; // @[IOManager.scala 123:13]
  wire  _GEN_81 = _GEN_79 & _GEN_80; // @[IOManager.scala 123:13]
  wire  _GEN_82 = ~_T_41; // @[IOManager.scala 139:13]
  wire  _GEN_83 = _T_38 & _GEN_82; // @[IOManager.scala 139:13]
  wire  _GEN_84 = ~_T_44; // @[IOManager.scala 139:13]
  wire  _GEN_85 = _GEN_83 & _GEN_84; // @[IOManager.scala 139:13]
  assign io_core_if__rdata = _T ? io_ram_rdata : _GEN_2; // @[IOManager.scala 66:7 IOManager.scala 74:16 IOManager.scala 74:16 IOManager.scala 74:16]
  assign io_core_if__ok = _T_38 ? _GEN_64 : _GEN_5; // @[IOManager.scala 66:7 IOManager.scala 75:13 IOManager.scala 75:13 IOManager.scala 75:13 IOManager.scala 133:14 IOManager.scala 137:14]
  assign io_core_mem_rdata = _T_3 ? io_ram_rdata : _GEN_8; // @[IOManager.scala 65:7 IOManager.scala 74:16 IOManager.scala 74:16 IOManager.scala 74:16]
  assign io_core_mem_ok = _T_18 ? _GEN_37 : _GEN_11; // @[IOManager.scala 65:7 IOManager.scala 75:13 IOManager.scala 75:13 IOManager.scala 75:13 IOManager.scala 103:16 IOManager.scala 106:16 IOManager.scala 117:16 IOManager.scala 120:16]
  assign io_ram_addr = _T_38 ? _GEN_61 : _GEN_45; // @[IOManager.scala 62:10 IOManager.scala 79:17 IOManager.scala 79:17]
  assign io_ram_mode = _T_38 ? _GEN_60 : _GEN_44; // @[IOManager.scala 62:10 IOManager.scala 78:17 IOManager.scala 78:17]
  assign io_ram_wdata = _T_38 ? _GEN_62 : _GEN_46; // @[IOManager.scala 62:10 IOManager.scala 80:18 IOManager.scala 80:18]
  assign io_flash_addr = _T_38 ? _GEN_66 : _GEN_50; // @[IOManager.scala 63:12 IOManager.scala 79:17 IOManager.scala 79:17]
  assign io_flash_mode = _T_38 ? _GEN_65 : _GEN_49; // @[IOManager.scala 63:12 IOManager.scala 78:17 IOManager.scala 78:17]
  assign io_flash_wdata = _T_38 ? _GEN_67 : _GEN_51; // @[IOManager.scala 63:12 IOManager.scala 80:18 IOManager.scala 80:18]
  assign io_serial_addr = _T_18 ? _GEN_42 : 32'h0; // @[IOManager.scala 64:13 IOManager.scala 79:17]
  assign io_serial_mode = _T_18 ? _GEN_41 : 4'h0; // @[IOManager.scala 64:13 IOManager.scala 78:17]
  assign io_serial_wdata = _T_18 ? _GEN_43 : 32'h0; // @[IOManager.scala 64:13 IOManager.scala 80:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ifWait = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  memWait = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ifWait <= 2'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        ifWait <= 2'h1;
      end else if (_T_44) begin
        ifWait <= 2'h2;
      end else if (!(_T_10)) begin
        ifWait <= 2'h0;
      end
    end else if (!(_T_10)) begin
      ifWait <= 2'h0;
    end
    if (reset) begin
      memWait <= 2'h0;
    end else if (_T_18) begin
      if (_T_21) begin
        if (io_core_mem_mode[3]) begin
          memWait <= 2'h0;
        end else begin
          memWait <= 2'h1;
        end
      end else if (_T_25) begin
        if (flashFree) begin
          memWait <= 2'h2;
        end else if (!(_T_14)) begin
          memWait <= 2'h0;
        end
      end else if (_T_28) begin
        if (io_core_mem_mode[3]) begin
          memWait <= 2'h0;
        end else begin
          memWait <= 2'h3;
        end
      end else if (!(_T_14)) begin
        memWait <= 2'h0;
      end
    end else if (!(_T_14)) begin
      memWait <= 2'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_81 & _T_31) begin
          $fwrite(32'h80000002,"[IO] MEM access invalid address: %x\n",io_core_mem_addr); // @[IOManager.scala 123:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_85 & _T_31) begin
          $fwrite(32'h80000002,"[IO] IF access invalid address: %x\n",io_core_if__addr); // @[IOManager.scala 139:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ChiselTop(
  input         clock,
  input         reset,
  output [31:0] io_ram_addr,
  output [3:0]  io_ram_mode,
  output [31:0] io_ram_wdata,
  input  [31:0] io_ram_rdata,
  input         io_ram_ok,
  output [31:0] io_flash_addr,
  output [3:0]  io_flash_mode,
  output [31:0] io_flash_wdata,
  input  [31:0] io_flash_rdata,
  input         io_flash_ok,
  output [31:0] io_serial_addr,
  output [3:0]  io_serial_mode,
  output [31:0] io_serial_wdata,
  input  [31:0] io_serial_rdata,
  input         io_serial_ok,
  output [31:0] io_debug_idex_aluOp_rd1,
  output [31:0] io_debug_idex_aluOp_rd2,
  output [4:0]  io_debug_idex_aluOp_opt,
  output [4:0]  io_debug_idex_wrRegOp_addr,
  output [31:0] io_debug_idex_wrRegOp_data,
  output        io_debug_idex_wrRegOp_rdy,
  output        io_debug_idex_wrCSROp_valid,
  output [11:0] io_debug_idex_wrCSROp_addr,
  output [31:0] io_debug_idex_wrCSROp_data,
  output [31:0] io_debug_idex_store_data,
  output        io_debug_idex_excep_valid,
  output [31:0] io_debug_idex_excep_code,
  output [31:0] io_debug_idex_excep_value,
  output [31:0] io_debug_idex_excep_pc,
  output        io_debug_idex_excep_valid_inst,
  output [31:0] io_debug_ifpc,
  output [31:0] io_debug_reg_0,
  output [31:0] io_debug_reg_1,
  output [31:0] io_debug_reg_2,
  output [31:0] io_debug_reg_3,
  output [31:0] io_debug_reg_4,
  output [31:0] io_debug_reg_5,
  output [31:0] io_debug_reg_6,
  output [31:0] io_debug_reg_7,
  output [31:0] io_debug_reg_8,
  output [31:0] io_debug_reg_9,
  output [31:0] io_debug_reg_10,
  output [31:0] io_debug_reg_11,
  output [31:0] io_debug_reg_12,
  output [31:0] io_debug_reg_13,
  output [31:0] io_debug_reg_14,
  output [31:0] io_debug_reg_15,
  output [31:0] io_debug_reg_16,
  output [31:0] io_debug_reg_17,
  output [31:0] io_debug_reg_18,
  output [31:0] io_debug_reg_19,
  output [31:0] io_debug_reg_20,
  output [31:0] io_debug_reg_21,
  output [31:0] io_debug_reg_22,
  output [31:0] io_debug_reg_23,
  output [31:0] io_debug_reg_24,
  output [31:0] io_debug_reg_25,
  output [31:0] io_debug_reg_26,
  output [31:0] io_debug_reg_27,
  output [31:0] io_debug_reg_28,
  output [31:0] io_debug_reg_29,
  output [31:0] io_debug_reg_30,
  output [31:0] io_debug_reg_31,
  output        io_debug_finish_pc_valid,
  output [31:0] io_debug_finish_pc_bits
);
  wire  core_clock; // @[Main.scala 16:23]
  wire  core_reset; // @[Main.scala 16:23]
  wire [31:0] core_io_dev_if__addr; // @[Main.scala 16:23]
  wire [3:0] core_io_dev_if__mode; // @[Main.scala 16:23]
  wire [31:0] core_io_dev_if__rdata; // @[Main.scala 16:23]
  wire  core_io_dev_if__ok; // @[Main.scala 16:23]
  wire [31:0] core_io_dev_mem_addr; // @[Main.scala 16:23]
  wire [3:0] core_io_dev_mem_mode; // @[Main.scala 16:23]
  wire [31:0] core_io_dev_mem_wdata; // @[Main.scala 16:23]
  wire [31:0] core_io_dev_mem_rdata; // @[Main.scala 16:23]
  wire  core_io_dev_mem_ok; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_aluOp_rd1; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_aluOp_rd2; // @[Main.scala 16:23]
  wire [4:0] core_io_debug_idex_aluOp_opt; // @[Main.scala 16:23]
  wire [4:0] core_io_debug_idex_wrRegOp_addr; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_wrRegOp_data; // @[Main.scala 16:23]
  wire  core_io_debug_idex_wrRegOp_rdy; // @[Main.scala 16:23]
  wire  core_io_debug_idex_wrCSROp_valid; // @[Main.scala 16:23]
  wire [11:0] core_io_debug_idex_wrCSROp_addr; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_wrCSROp_data; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_store_data; // @[Main.scala 16:23]
  wire  core_io_debug_idex_excep_valid; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_excep_code; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_excep_value; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_idex_excep_pc; // @[Main.scala 16:23]
  wire  core_io_debug_idex_excep_valid_inst; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_ifpc; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_0; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_1; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_2; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_3; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_4; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_5; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_6; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_7; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_8; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_9; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_10; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_11; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_12; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_13; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_14; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_15; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_16; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_17; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_18; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_19; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_20; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_21; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_22; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_23; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_24; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_25; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_26; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_27; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_28; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_29; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_30; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_reg_31; // @[Main.scala 16:23]
  wire  core_io_debug_finish_pc_valid; // @[Main.scala 16:23]
  wire [31:0] core_io_debug_finish_pc_bits; // @[Main.scala 16:23]
  wire  ioCtrl_clock; // @[Main.scala 17:23]
  wire  ioCtrl_reset; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_core_if__addr; // @[Main.scala 17:23]
  wire [3:0] ioCtrl_io_core_if__mode; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_core_if__rdata; // @[Main.scala 17:23]
  wire  ioCtrl_io_core_if__ok; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_core_mem_addr; // @[Main.scala 17:23]
  wire [3:0] ioCtrl_io_core_mem_mode; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_core_mem_wdata; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_core_mem_rdata; // @[Main.scala 17:23]
  wire  ioCtrl_io_core_mem_ok; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_ram_addr; // @[Main.scala 17:23]
  wire [3:0] ioCtrl_io_ram_mode; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_ram_wdata; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_ram_rdata; // @[Main.scala 17:23]
  wire  ioCtrl_io_ram_ok; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_flash_addr; // @[Main.scala 17:23]
  wire [3:0] ioCtrl_io_flash_mode; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_flash_wdata; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_flash_rdata; // @[Main.scala 17:23]
  wire  ioCtrl_io_flash_ok; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_serial_addr; // @[Main.scala 17:23]
  wire [3:0] ioCtrl_io_serial_mode; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_serial_wdata; // @[Main.scala 17:23]
  wire [31:0] ioCtrl_io_serial_rdata; // @[Main.scala 17:23]
  wire  ioCtrl_io_serial_ok; // @[Main.scala 17:23]
  Core core ( // @[Main.scala 16:23]
    .clock(core_clock),
    .reset(core_reset),
    .io_dev_if__addr(core_io_dev_if__addr),
    .io_dev_if__mode(core_io_dev_if__mode),
    .io_dev_if__rdata(core_io_dev_if__rdata),
    .io_dev_if__ok(core_io_dev_if__ok),
    .io_dev_mem_addr(core_io_dev_mem_addr),
    .io_dev_mem_mode(core_io_dev_mem_mode),
    .io_dev_mem_wdata(core_io_dev_mem_wdata),
    .io_dev_mem_rdata(core_io_dev_mem_rdata),
    .io_dev_mem_ok(core_io_dev_mem_ok),
    .io_debug_idex_aluOp_rd1(core_io_debug_idex_aluOp_rd1),
    .io_debug_idex_aluOp_rd2(core_io_debug_idex_aluOp_rd2),
    .io_debug_idex_aluOp_opt(core_io_debug_idex_aluOp_opt),
    .io_debug_idex_wrRegOp_addr(core_io_debug_idex_wrRegOp_addr),
    .io_debug_idex_wrRegOp_data(core_io_debug_idex_wrRegOp_data),
    .io_debug_idex_wrRegOp_rdy(core_io_debug_idex_wrRegOp_rdy),
    .io_debug_idex_wrCSROp_valid(core_io_debug_idex_wrCSROp_valid),
    .io_debug_idex_wrCSROp_addr(core_io_debug_idex_wrCSROp_addr),
    .io_debug_idex_wrCSROp_data(core_io_debug_idex_wrCSROp_data),
    .io_debug_idex_store_data(core_io_debug_idex_store_data),
    .io_debug_idex_excep_valid(core_io_debug_idex_excep_valid),
    .io_debug_idex_excep_code(core_io_debug_idex_excep_code),
    .io_debug_idex_excep_value(core_io_debug_idex_excep_value),
    .io_debug_idex_excep_pc(core_io_debug_idex_excep_pc),
    .io_debug_idex_excep_valid_inst(core_io_debug_idex_excep_valid_inst),
    .io_debug_ifpc(core_io_debug_ifpc),
    .io_debug_reg_0(core_io_debug_reg_0),
    .io_debug_reg_1(core_io_debug_reg_1),
    .io_debug_reg_2(core_io_debug_reg_2),
    .io_debug_reg_3(core_io_debug_reg_3),
    .io_debug_reg_4(core_io_debug_reg_4),
    .io_debug_reg_5(core_io_debug_reg_5),
    .io_debug_reg_6(core_io_debug_reg_6),
    .io_debug_reg_7(core_io_debug_reg_7),
    .io_debug_reg_8(core_io_debug_reg_8),
    .io_debug_reg_9(core_io_debug_reg_9),
    .io_debug_reg_10(core_io_debug_reg_10),
    .io_debug_reg_11(core_io_debug_reg_11),
    .io_debug_reg_12(core_io_debug_reg_12),
    .io_debug_reg_13(core_io_debug_reg_13),
    .io_debug_reg_14(core_io_debug_reg_14),
    .io_debug_reg_15(core_io_debug_reg_15),
    .io_debug_reg_16(core_io_debug_reg_16),
    .io_debug_reg_17(core_io_debug_reg_17),
    .io_debug_reg_18(core_io_debug_reg_18),
    .io_debug_reg_19(core_io_debug_reg_19),
    .io_debug_reg_20(core_io_debug_reg_20),
    .io_debug_reg_21(core_io_debug_reg_21),
    .io_debug_reg_22(core_io_debug_reg_22),
    .io_debug_reg_23(core_io_debug_reg_23),
    .io_debug_reg_24(core_io_debug_reg_24),
    .io_debug_reg_25(core_io_debug_reg_25),
    .io_debug_reg_26(core_io_debug_reg_26),
    .io_debug_reg_27(core_io_debug_reg_27),
    .io_debug_reg_28(core_io_debug_reg_28),
    .io_debug_reg_29(core_io_debug_reg_29),
    .io_debug_reg_30(core_io_debug_reg_30),
    .io_debug_reg_31(core_io_debug_reg_31),
    .io_debug_finish_pc_valid(core_io_debug_finish_pc_valid),
    .io_debug_finish_pc_bits(core_io_debug_finish_pc_bits)
  );
  IOManager ioCtrl ( // @[Main.scala 17:23]
    .clock(ioCtrl_clock),
    .reset(ioCtrl_reset),
    .io_core_if__addr(ioCtrl_io_core_if__addr),
    .io_core_if__mode(ioCtrl_io_core_if__mode),
    .io_core_if__rdata(ioCtrl_io_core_if__rdata),
    .io_core_if__ok(ioCtrl_io_core_if__ok),
    .io_core_mem_addr(ioCtrl_io_core_mem_addr),
    .io_core_mem_mode(ioCtrl_io_core_mem_mode),
    .io_core_mem_wdata(ioCtrl_io_core_mem_wdata),
    .io_core_mem_rdata(ioCtrl_io_core_mem_rdata),
    .io_core_mem_ok(ioCtrl_io_core_mem_ok),
    .io_ram_addr(ioCtrl_io_ram_addr),
    .io_ram_mode(ioCtrl_io_ram_mode),
    .io_ram_wdata(ioCtrl_io_ram_wdata),
    .io_ram_rdata(ioCtrl_io_ram_rdata),
    .io_ram_ok(ioCtrl_io_ram_ok),
    .io_flash_addr(ioCtrl_io_flash_addr),
    .io_flash_mode(ioCtrl_io_flash_mode),
    .io_flash_wdata(ioCtrl_io_flash_wdata),
    .io_flash_rdata(ioCtrl_io_flash_rdata),
    .io_flash_ok(ioCtrl_io_flash_ok),
    .io_serial_addr(ioCtrl_io_serial_addr),
    .io_serial_mode(ioCtrl_io_serial_mode),
    .io_serial_wdata(ioCtrl_io_serial_wdata),
    .io_serial_rdata(ioCtrl_io_serial_rdata),
    .io_serial_ok(ioCtrl_io_serial_ok)
  );
  assign io_ram_addr = ioCtrl_io_ram_addr; // @[Main.scala 21:15]
  assign io_ram_mode = ioCtrl_io_ram_mode; // @[Main.scala 21:15]
  assign io_ram_wdata = ioCtrl_io_ram_wdata; // @[Main.scala 21:15]
  assign io_flash_addr = ioCtrl_io_flash_addr; // @[Main.scala 22:15]
  assign io_flash_mode = ioCtrl_io_flash_mode; // @[Main.scala 22:15]
  assign io_flash_wdata = ioCtrl_io_flash_wdata; // @[Main.scala 22:15]
  assign io_serial_addr = ioCtrl_io_serial_addr; // @[Main.scala 23:15]
  assign io_serial_mode = ioCtrl_io_serial_mode; // @[Main.scala 23:15]
  assign io_serial_wdata = ioCtrl_io_serial_wdata; // @[Main.scala 23:15]
  assign io_debug_idex_aluOp_rd1 = core_io_debug_idex_aluOp_rd1; // @[Main.scala 20:17]
  assign io_debug_idex_aluOp_rd2 = core_io_debug_idex_aluOp_rd2; // @[Main.scala 20:17]
  assign io_debug_idex_aluOp_opt = core_io_debug_idex_aluOp_opt; // @[Main.scala 20:17]
  assign io_debug_idex_wrRegOp_addr = core_io_debug_idex_wrRegOp_addr; // @[Main.scala 20:17]
  assign io_debug_idex_wrRegOp_data = core_io_debug_idex_wrRegOp_data; // @[Main.scala 20:17]
  assign io_debug_idex_wrRegOp_rdy = core_io_debug_idex_wrRegOp_rdy; // @[Main.scala 20:17]
  assign io_debug_idex_wrCSROp_valid = core_io_debug_idex_wrCSROp_valid; // @[Main.scala 20:17]
  assign io_debug_idex_wrCSROp_addr = core_io_debug_idex_wrCSROp_addr; // @[Main.scala 20:17]
  assign io_debug_idex_wrCSROp_data = core_io_debug_idex_wrCSROp_data; // @[Main.scala 20:17]
  assign io_debug_idex_store_data = core_io_debug_idex_store_data; // @[Main.scala 20:17]
  assign io_debug_idex_excep_valid = core_io_debug_idex_excep_valid; // @[Main.scala 20:17]
  assign io_debug_idex_excep_code = core_io_debug_idex_excep_code; // @[Main.scala 20:17]
  assign io_debug_idex_excep_value = core_io_debug_idex_excep_value; // @[Main.scala 20:17]
  assign io_debug_idex_excep_pc = core_io_debug_idex_excep_pc; // @[Main.scala 20:17]
  assign io_debug_idex_excep_valid_inst = core_io_debug_idex_excep_valid_inst; // @[Main.scala 20:17]
  assign io_debug_ifpc = core_io_debug_ifpc; // @[Main.scala 20:17]
  assign io_debug_reg_0 = core_io_debug_reg_0; // @[Main.scala 20:17]
  assign io_debug_reg_1 = core_io_debug_reg_1; // @[Main.scala 20:17]
  assign io_debug_reg_2 = core_io_debug_reg_2; // @[Main.scala 20:17]
  assign io_debug_reg_3 = core_io_debug_reg_3; // @[Main.scala 20:17]
  assign io_debug_reg_4 = core_io_debug_reg_4; // @[Main.scala 20:17]
  assign io_debug_reg_5 = core_io_debug_reg_5; // @[Main.scala 20:17]
  assign io_debug_reg_6 = core_io_debug_reg_6; // @[Main.scala 20:17]
  assign io_debug_reg_7 = core_io_debug_reg_7; // @[Main.scala 20:17]
  assign io_debug_reg_8 = core_io_debug_reg_8; // @[Main.scala 20:17]
  assign io_debug_reg_9 = core_io_debug_reg_9; // @[Main.scala 20:17]
  assign io_debug_reg_10 = core_io_debug_reg_10; // @[Main.scala 20:17]
  assign io_debug_reg_11 = core_io_debug_reg_11; // @[Main.scala 20:17]
  assign io_debug_reg_12 = core_io_debug_reg_12; // @[Main.scala 20:17]
  assign io_debug_reg_13 = core_io_debug_reg_13; // @[Main.scala 20:17]
  assign io_debug_reg_14 = core_io_debug_reg_14; // @[Main.scala 20:17]
  assign io_debug_reg_15 = core_io_debug_reg_15; // @[Main.scala 20:17]
  assign io_debug_reg_16 = core_io_debug_reg_16; // @[Main.scala 20:17]
  assign io_debug_reg_17 = core_io_debug_reg_17; // @[Main.scala 20:17]
  assign io_debug_reg_18 = core_io_debug_reg_18; // @[Main.scala 20:17]
  assign io_debug_reg_19 = core_io_debug_reg_19; // @[Main.scala 20:17]
  assign io_debug_reg_20 = core_io_debug_reg_20; // @[Main.scala 20:17]
  assign io_debug_reg_21 = core_io_debug_reg_21; // @[Main.scala 20:17]
  assign io_debug_reg_22 = core_io_debug_reg_22; // @[Main.scala 20:17]
  assign io_debug_reg_23 = core_io_debug_reg_23; // @[Main.scala 20:17]
  assign io_debug_reg_24 = core_io_debug_reg_24; // @[Main.scala 20:17]
  assign io_debug_reg_25 = core_io_debug_reg_25; // @[Main.scala 20:17]
  assign io_debug_reg_26 = core_io_debug_reg_26; // @[Main.scala 20:17]
  assign io_debug_reg_27 = core_io_debug_reg_27; // @[Main.scala 20:17]
  assign io_debug_reg_28 = core_io_debug_reg_28; // @[Main.scala 20:17]
  assign io_debug_reg_29 = core_io_debug_reg_29; // @[Main.scala 20:17]
  assign io_debug_reg_30 = core_io_debug_reg_30; // @[Main.scala 20:17]
  assign io_debug_reg_31 = core_io_debug_reg_31; // @[Main.scala 20:17]
  assign io_debug_finish_pc_valid = core_io_debug_finish_pc_valid; // @[Main.scala 20:17]
  assign io_debug_finish_pc_bits = core_io_debug_finish_pc_bits; // @[Main.scala 20:17]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_dev_if__rdata = ioCtrl_io_core_if__rdata; // @[Main.scala 19:15]
  assign core_io_dev_if__ok = ioCtrl_io_core_if__ok; // @[Main.scala 19:15]
  assign core_io_dev_mem_rdata = ioCtrl_io_core_mem_rdata; // @[Main.scala 19:15]
  assign core_io_dev_mem_ok = ioCtrl_io_core_mem_ok; // @[Main.scala 19:15]
  assign ioCtrl_clock = clock;
  assign ioCtrl_reset = reset;
  assign ioCtrl_io_core_if__addr = core_io_dev_if__addr; // @[Main.scala 19:15]
  assign ioCtrl_io_core_if__mode = core_io_dev_if__mode; // @[Main.scala 19:15]
  assign ioCtrl_io_core_mem_addr = core_io_dev_mem_addr; // @[Main.scala 19:15]
  assign ioCtrl_io_core_mem_mode = core_io_dev_mem_mode; // @[Main.scala 19:15]
  assign ioCtrl_io_core_mem_wdata = core_io_dev_mem_wdata; // @[Main.scala 19:15]
  assign ioCtrl_io_ram_rdata = io_ram_rdata; // @[Main.scala 21:15]
  assign ioCtrl_io_ram_ok = io_ram_ok; // @[Main.scala 21:15]
  assign ioCtrl_io_flash_rdata = io_flash_rdata; // @[Main.scala 22:15]
  assign ioCtrl_io_flash_ok = io_flash_ok; // @[Main.scala 22:15]
  assign ioCtrl_io_serial_rdata = io_serial_rdata; // @[Main.scala 23:15]
  assign ioCtrl_io_serial_ok = io_serial_ok; // @[Main.scala 23:15]
endmodule
